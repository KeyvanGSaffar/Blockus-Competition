library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std.All;

-------------------------------
---- Uncomment the following library declaration if instantiating
entity program_coding is
    Port ( datain :in std_logic_vector (117 downto 0);
				  data_coded :  out std_logic_vector(31 downto 0)
);
end program_coding;
-------------------------------------
architecture Gate_level of program_coding is

		type MATRIX is array(5 downto 0) of std_logic_vector(17 downto 0);

		signal X_black_before,Y_black_before : unsigned(4 downto 0);
		signal X_black,Y_black : unsigned (7 downto 0);
		signal format : unsigned (7 downto 0);
		signal rotate : unsigned (7 downto 0);
		
		type MAT_ATTACHED is array(7 downto 0) of std_logic_vector(107 downto 0);
		signal sampler : std_logic_vector(107 downto 0) := (others=>'0');
--		signal a,b,c,d,e,f,g,h,i,j,k,l,m,n,o,p,q	:	MAT_ATTACHED;


--
--		constant a_0 :MATRIX :=( "000000000000000000","000000000000000000","000011010011000000","000010100010000000","000011010011000000","000000000000000000");
--		constant a_1 :MATRIX :=(	"000000000000000000","000000000000000000","000000011010011000","000000010100010000","000000011010011000","000000000000000000");
--		constant a_2 :MATRIX :=( "000000000000000000","000011010011000000","000010100010000000","000011010011000000","000000000000000000","000000000000000000");
--		constant a_3 :MATRIX :=( "000000000000000000","000000011010011000","000000010100010000","000000011010011000","000000000000000000","000000000000000000");
--		constant a_4 :MATRIX :=( "000000000000000000","000011010011000000","000010100010000000","000011010011000000","000000000000000000","000000000000000000");
--		constant a_5 :MATRIX :=( "000000000000000000","000000011010011000","000000010100010000","000000011010011000","000000000000000000","000000000000000000");
--		constant a_6 :MATRIX :=( "000000000000000000","000000000000000000","000011010011000000","000010100010000000","000011010011000000","000000000000000000");
--		constant a_7 :MATRIX :=( "000000000000000000","000000000000000000","000000011010011000","000000010100010000","000000011010011000","000000000000000000");
--		constant b_0 :MATRIX :=( "000000000000000000","000000000000000000","000011010011000000","000010100010000000","000010001010000000","000011010011000000");
--		constant b_1 :MATRIX :=( "000000000000000000","000000000000000000","000000011010011000","000000010100010000","000000010001010000","000000011010011000");
--		constant b_2 :MATRIX :=( "000011010011000000","000010001010000000","000010100010000000","000011010011000000","000000000000000000","000000000000000000");
--		constant b_3 :MATRIX :=( "000000011010011000","000000010001010000","000000010100010000","000000011010011000","000000000000000000","000000000000000000");
--		constant b_4 :MATRIX :=( "000000000000000000","011010010011000000","010001100010000000","011010010011000000","000000000000000000","000000000000000000");
--		constant b_5 :MATRIX :=( "000000000000000000","000000011010010011","000000010100001010","000000011010010011","000000000000000000","000000000000000000");
--		constant b_6 :MATRIX :=( "000000000000000000","000000000000000000","011010010011000000","010001100010000000","011010010011000000","000000000000000000");
--		constant b_7 :MATRIX :=( "000000000000000000","000000000000000000","000000011010010011","000000010100001010","000000011010010011","000000000000000000");
--		constant c_0 :MATRIX :=( "000000000000000000","000011010011000000","000010001010000000","000010100010000000","000010001010000000","000011010011000000");
--		constant c_1 :MATRIX :=( "000000000000000000","000000011010011000","000000010001010000","000000010100010000","000000010001010000","000000011010011000");
--		constant c_2 :MATRIX :=( "000011010011000000","000010001010000000","000010100010000000","000010001010000000","000011010011000000","000000000000000000");
--		constant c_3 :MATRIX :=( "000000011010011000","000000010001010000","000000010100010000","000000010001010000","000000011010011000","000000000000000000");
--		constant c_4 :MATRIX :=( "000000000000000000","011010010010011000","010001100001010000","011010010010011000","000000000000000000","000000000000000000");
--		constant c_5 :MATRIX :=( "000000000000000000","000011010010010011","000010001100001010","000011010010010011","000000000000000000","000000000000000000");
--		constant c_6 :MATRIX :=( "000000000000000000","000000000000000000","011010010010011000","010001100001010000","011010010010011000","000000000000000000");
--		constant c_7 :MATRIX :=( "000000000000000000","000000000000000000","000011010010010011","000010001100001010","000011010010010011","000000000000000000");
--		constant d_0 :MATRIX :=( "000000000000000000","000011010011000000","000010001010011000","000010100001010000","000011010010011000","000000000000000000");
--		constant d_1 :MATRIX :=( "000000000000000000","000000011010011000","000011010001010000","000010001100010000","000011010010011000","000000000000000000");
--		constant d_2 :MATRIX :=( "000000000000000000","000011010010011000","000010100001010000","000010001010011000","000011010011000000","000000000000000000");
--		constant d_3 :MATRIX :=( "000000000000000000","000011010010011000","000010001100010000","000011010001010000","000000011010011000","000000000000000000");
--		constant d_4 :MATRIX :=( "000000000000000000","000011010010011000","000010100001010000","000010001010011000","000011010011000000","000000000000000000");
--		constant d_5 :MATRIX :=( "000000000000000000","000011010010011000","000010001100010000","000011010001010000","000000011010011000","000000000000000000");
--		constant d_6 :MATRIX :=( "000000000000000000","000011010011000000","000010001010011000","000010100001010000","000011010010011000","000000000000000000");
--		constant d_7 :MATRIX :=( "000000000000000000","000000011010011000","000011010001010000","000010001100010000","000011010010011000","000000000000000000");
--		constant e_0 :MATRIX :=( "000000000000000000","000011010011000000","000010001010000000","011010100010000000","010001001010000000","011010010011000000");
--		constant e_1 :MATRIX :=( "000000000000000000","000000011010011000","000000010001010000","000000010100010011","000000010001001010","000000011010010011");
--		constant e_2 :MATRIX :=( "011010010011000000","010001001010000000","011010100010000000","000010001010000000","000011010011000000","000000000000000000");
--		constant e_3 :MATRIX :=( "000000011010010011","000000010001001010","000000010100010011","000000010001010000","000000011010011000","000000000000000000");
--		constant e_4 :MATRIX :=( "011010011000000000","010001010010011000","010001100001010000","011010010010011000","000000000000000000","000000000000000000");
--		constant e_5 :MATRIX :=( "000000000011010011","000011010010001010","000010001100001010","000011010010010011","000000000000000000","000000000000000000");
--		constant e_6 :MATRIX :=( "000000000000000000","000000000000000000","011010010010011000","010001100001010000","010001010010011000","011010011000000000");
--		constant e_7 :MATRIX :=( "000000000000000000","000000000000000000","000011010010010011","000010001100001010","000011010010001010","000000000011010011");
--		constant f_0 :MATRIX :=( "000000000000000000","000011010011000000","000010001010011000","000010100001010000","000010001010011000","000011010011000000");
--		constant f_1 :MATRIX :=( "000000000000000000","000000011010011000","000011010001010000","000010001100010000","000011010001010000","000000011010011000");
--		constant f_2 :MATRIX :=( "000011010011000000","000010001010011000","000010100001010000","000010001010011000","000011010011000000","000000000000000000");
--		constant f_3 :MATRIX :=( "000000011010011000","000011010001010000","000010001100010000","000011010001010000","000000011010011000","000000000000000000");
--		constant f_4 :MATRIX :=( "000000000000000000","011010010010011000","010001100001010000","011010001010011000","000011010011000000","000000000000000000");
--		constant f_5 :MATRIX :=( "000000000000000000","000011010010010011","000010001100001010","000011010001010011","000000011010011000","000000000000000000");
--		constant f_6 :MATRIX :=( "000000000000000000","000011010011000000","011010001010011000","010001100001010000","011010010010011000","000000000000000000");
--		constant f_7 :MATRIX :=( "000000000000000000","000000011010011000","000011010001010011","000010001100001010","000011010010010011","000000000000000000");
--		constant g_0 :MATRIX :=( "000000000000000000","000000000000000000","000011010010011000","000010100001010000","000010001001010000","000011010010011000");
--		constant g_1 :MATRIX :=( "000000000000000000","000000000000000000","000011010010011000","000010001100010000","000010001001010000","000011010010011000");
--		constant g_2 :MATRIX :=( "000011010010011000","000010001001010000","000010100001010000","000011010010011000","000000000000000000","000000000000000000");
--		constant g_3 :MATRIX :=( "000011010010011000","000010001001010000","000010001100010000","000011010010011000","000000000000000000","000000000000000000");
--		constant g_4 :MATRIX :=( "000000000000000000","011010010011000000","010001100010000000","010001001010000000","011010010011000000","000000000000000000");
--		constant g_5 :MATRIX :=( "000000000000000000","000000011010010011","000000010100001010","000000010001001010","000000011010010011","000000000000000000");
--		constant g_6 :MATRIX :=( "000000000000000000","011010010011000000","010001001010000000","010001100010000000","011010010011000000","000000000000000000");
--		constant g_7 :MATRIX :=( "000000000000000000","000000011010010011","000000010001001010","000000010100001010","000000011010010011","000000000000000000");
--		constant h_0 :MATRIX :=( "000000000000000000","000000000000000000","011010010011000000","010001100010011000","011010001001010000","000011010010011000");
--		constant h_1 :MATRIX :=( "000000000000000000","000000000000000000","000000011010010011","000011010100001010","000010001001010011","000011010010011000");
--		constant h_2 :MATRIX :=( "000011010010011000","011010001001010000","010001100010011000","011010010011000000","000000000000000000","000000000000000000");
--		constant h_3 :MATRIX :=( "000011010010011000","000010001001010011","000011010100001010","000000011010010011","000000000000000000","000000000000000000");
--		constant h_4 :MATRIX :=( "000011010011000000","011010001010000000","010001100010000000","010001010011000000","011010011000000000","000000000000000000");
--		constant h_5 :MATRIX :=( "000000011010011000","000000010001010011","000000010100001010","000000011010001010","000000000011010011","000000000000000000");
--		constant h_6 :MATRIX :=( "000000000000000000","011010011000000000","010001010011000000","010001100010000000","011010001010000000","000011010011000000");
--		constant h_7 :MATRIX :=( "000000000000000000","000000000011010011","000000011010001010","000000010100001010","000000010001010011","000000011010011000");
--		constant i_0 :MATRIX :=( "000011010011000000","000010001010000000","011010001010000000","010001100010000000","010001010011000000","011010011000000000");
--		constant i_1 :MATRIX :=( "000000011010011000","000000010001010000","000000010001010011","000000010100001010","000000011010001010","000000000011010011");
--		constant i_2 :MATRIX :=( "011010011000000000","010001010011000000","010001100010000000","011010001010000000","000010001010000000","000011010011000000");
--		constant i_3 :MATRIX :=( "000000000011010011","000000011010001010","000000010100001010","000000010001010011","000000010001010000","000000011010011000");
--		constant i_4 :MATRIX :=( "011010010011000000","010001001010010011","011010100001001010","000011010010010011","000000000000000000","000000000000000000");
--		constant i_5 :MATRIX :=( "000000011010010011","011010010001001010","010001001100010011","011010010010011000","000000000000000000","000000000000000000");
--		constant i_6 :MATRIX :=( "000000000000000000","000000000000000000","000011010010010011","011010100001001010","010001001010010011","011010010011000000");
--		constant i_7 :MATRIX :=( "000000000000000000","000000000000000000","011010010010011000","010001001100010011","011010010001001010","000000011010010011");
--		constant j_0 :MATRIX :=( "000000000000000000","000011010011000000","011010001010000000","010001100010000000","010001001010000000","011010010011000000");
--		constant j_1 :MATRIX :=( "000000000000000000","000000011010011000","000000010001010011","000000010100001010","000000010001001010","000000011010010011");
--		constant j_2 :MATRIX :=( "011010010011000000","010001001010000000","010001100010000000","011010001010000000","000011010011000000","000000000000000000");
--		constant j_3 :MATRIX :=( "000000011010010011","000000010001001010","000000010100001010","000000010001010011","000000011010011000","000000000000000000");
--		constant j_4 :MATRIX :=( "011010010011000000","010001001010011000","010001100001010000","011010010010011000","000000000000000000","000000000000000000");
--		constant j_5 :MATRIX :=( "000000011010010011","000011010001001010","000010001100001010","000011010010010011","000000000000000000","000000000000000000");
--		constant j_6 :MATRIX :=( "000000000000000000","000000000000000000","011010010010011000","010001100001010000","010001001010011000","011010010011000000");
--		constant j_7 :MATRIX :=( "000000000000000000","000000000000000000","000011010010010011","000010001100001010","000011010001001010","000000011010010011");
--		constant k_0 :MATRIX :=( "000000000000000000","011010010011000000","010001001010000000","011010100010000000","010001001010000000","011010010011000000");
--		constant k_1 :MATRIX :=( "000000000000000000","000000011010010011","000000010001001010","000000010100010011","000000010001001010","000000011010010011");
--		constant k_2 :MATRIX :=( "011010010011000000","010001001010000000","011010100010000000","010001001010000000","011010010011000000","000000000000000000");
--		constant k_3 :MATRIX :=( "000000011010010011","000000010001001010","000000010100010011","000000010001001010","000000011010010011","000000000000000000");
--		constant k_4 :MATRIX :=( "011010011010011000","010001010001010000","010001100001010000","011010010010011000","000000000000000000","000000000000000000");
--		constant k_5 :MATRIX :=( "000011010011010011","000010001010001010","000010001100001010","000011010010010011","000000000000000000","000000000000000000");
--		constant k_6 :MATRIX :=( "000000000000000000","000000000000000000","011010010010011000","010001100001010000","010001010001010000","011010011010011000");
--		constant k_7 :MATRIX :=( "000000000000000000","000000000000000000","000011010010010011","000010001100001010","000010001010001010","000011010011010011");
--		constant l_0 :MATRIX :=( "000000000000000000","000011010011000000","000010001010000000","011010100010011000","010001001001010000","011010010010011000");
--		constant l_1 :MATRIX :=( "000000000000000000","000000011010011000","000000010001010000","000011010100010011","000010001001001010","000011010010010011");
--		constant l_2 :MATRIX :=( "011010010010011000","010001001001010000","011010100010011000","000010001010000000","000011010011000000","000000000000000000");
--		constant l_3 :MATRIX :=( "000011010010010011","000010001001001010","000011010100010011","000000010001010000","000000011010011000","000000000000000000");
--		constant l_4 :MATRIX :=( "011010011000000000","010001010010011000","010001100001010000","010001010010011000","011010011000000000","000000000000000000");
--		constant l_5 :MATRIX :=( "000000000011010011","000011010010001010","000010001100001010","000011010010001010","000000000011010011","000000000000000000");
--		constant l_6 :MATRIX :=( "000000000000000000","011010011000000000","010001010010011000","010001100001010000","010001010010011000","011010011000000000");
--		constant l_7 :MATRIX :=( "000000000000000000","000000000011010011","000011010010001010","000010001100001010","000011010010001010","000000000011010011");
--		constant m_0 :MATRIX :=( "000011010011000000","000010001010000000","000010001010010011","000010100001001010","000011010010010011","000000000000000000");
--		constant m_1 :MATRIX :=( "000000011010011000","000000010001010000","011010010001010000","010001001100010000","011010010010011000","000000000000000000");
--		constant m_2 :MATRIX :=( "000000000000000000","000011010010010011","000010100001001010","000010001010010011","000010001010000000","000011010011000000");
--		constant m_3 :MATRIX :=( "000000000000000000","011010010010011000","010001001100010000","011010010001010000","000000010001010000","000000011010011000");
--		constant m_4 :MATRIX :=( "000000000000000000","000011010010010011","000010100001001010","000010001010010011","000010001010000000","000011010011000000");
--		constant m_5 :MATRIX :=( "000000000000000000","011010010010011000","010001001100010000","011010010001010000","000000010001010000","000000011010011000");
--		constant m_6 :MATRIX :=( "000011010011000000","000010001010000000","000010001010010011","000010100001001010","000011010010010011","000000000000000000");
--		constant m_7 :MATRIX :=( "000000011010011000","000000010001010000","011010010001010000","010001001100010000","011010010010011000","000000000000000000");
--		constant n_0 :MATRIX :=( "000000000000000000","011010010011000000","010001001010011000","011010100001010000","000011010001010000","000000011010011000");
--		constant n_1 :MATRIX :=( "000000000000000000","000000011010010011","000011010001001010","000010001100010011","000010001010011000","000011010011000000");
--		constant n_2 :MATRIX :=( "000000011010011000","000011010001010000","011010100001010000","010001001010011000","011010010011000000","000000000000000000");
--		constant n_3 :MATRIX :=( "000011010011000000","000010001010011000","000010001100010011","000011010001001010","000000011010010011","000000000000000000");
--		constant n_4 :MATRIX :=( "000000011010011000","000011010001010000","011010100001010000","010001001010011000","011010010011000000","000000000000000000");
--		constant n_5 :MATRIX :=( "000011010011000000","000010001010011000","000010001100010011","000011010001001010","000000011010010011","000000000000000000");
--		constant n_6 :MATRIX :=( "000000000000000000","011010010011000000","010001001010011000","011010100001010000","000011010001010000","000000011010011000");
--		constant n_7 :MATRIX :=( "000000000000000000","000000011010010011","000011010001001010","000010001100010011","000010001010011000","000011010011000000");
--		constant o_0 :MATRIX :=( "000000000000000000","011010011000000000","010001010010011000","010001100001010000","011010010001010000","000000011010011000");
--		constant o_1 :MATRIX :=( "000000000000000000","000000000011010011","000011010010001010","000010001100001010","000010001010010011","000011010011000000");
--		constant o_2 :MATRIX :=( "000000011010011000","011010010001010000","010001100001010000","010001010010011000","011010011000000000","000000000000000000");
--		constant o_3 :MATRIX :=( "000011010011000000","000010001010010011","000010001100001010","000011010010001010","000000000011010011","000000000000000000");
--		constant o_4 :MATRIX :=( "000011010010011000","000010001001010000","011010100010011000","010001001010000000","011010010011000000","000000000000000000");
--		constant o_5 :MATRIX :=( "000011010010011000","000010001001010000","000011010100010011","000000010001001010","000000011010010011","000000000000000000");
--		constant o_6 :MATRIX :=( "000000000000000000","011010010011000000","010001001010000000","011010100010011000","000010001001010000","000011010010011000");
--		constant o_7 :MATRIX :=( "000000000000000000","000000011010010011","000000010001001010","000011010100010011","000010001001010000","000011010010011000");
--		constant p_0 :MATRIX :=( "000000000000000000","011010011000000000","010001010010011000","010001100001010000","011010001010011000","000011010011000000");
--		constant p_1 :MATRIX :=( "000000000000000000","000000000011010011","000011010010001010","000010001100001010","000011010001010011","000000011010011000");
--		constant p_2 :MATRIX :=( "000011010011000000","011010001010011000","010001100001010000","010001010010011000","011010011000000000","000000000000000000");
--		constant p_3 :MATRIX :=( "000000011010011000","000011010001010011","000010001100001010","000011010010001010","000000000011010011","000000000000000000");
--		constant p_4 :MATRIX :=( "000011010010011000","011010001001010000","010001100010011000","011010001010000000","000011010011000000","000000000000000000");
--		constant p_5 :MATRIX :=( "000011010010011000","000010001001010011","000011010100001010","000000010001010011","000000011010011000","000000000000000000");
--		constant p_6 :MATRIX :=( "000000000000000000","000011010011000000","011010001010000000","010001100010011000","011010001001010000","000011010010011000");
--		constant p_7 :MATRIX :=( "000000000000000000","000000011010011000","000000010001010011","000011010100001010","000010001001010011","000011010010011000");
--		constant q_0 :MATRIX :=( "000000000000000000","000011010011000000","011010001010011000","010001100001010000","011010001010011000","000011010011000000");
--		constant q_1 :MATRIX :=( "000000000000000000","000000011010011000","000011010001010011","000010001100001010","000011010001010011","000000011010011000");
--		constant q_2 :MATRIX :=( "000011010011000000","011010001010011000","010001100001010000","011010001010011000","000011010011000000","000000000000000000");
--		constant q_3 :MATRIX :=( "000000011010011000","000011010001010011","000010001100001010","000011010001010011","000000011010011000","000000000000000000");
--		constant q_4 :MATRIX :=( "000011010011000000","011010001010011000","010001100001010000","011010001010011000","000011010011000000","000000000000000000");
--		constant q_5 :MATRIX :=( "000000011010011000","000011010001010011","000010001100001010","000011010001010011","000000011010011000","000000000000000000");
--		constant q_6 :MATRIX :=( "000000000000000000","000011010011000000","011010001010011000","010001100001010000","011010001010011000","000011010011000000");
--		constant q_7 :MATRIX :=(	"000000000000000000","000000011010011000","000011010001010011","000010001100001010","000011010001010011","000000011010011000");
--
--

		constant a_0 :std_logic_vector(107 downto 0) :=( "000000000000000000000000000000000000000011010011000000000010100010000000000011010011000000000000000000000000");
		constant a_1 :std_logic_vector(107 downto 0) :=( "000000000000000000000000000000000000000000011010011000000000010100010000000000011010011000000000000000000000");
		constant a_2 :std_logic_vector(107 downto 0) :=( "000000000000000000000011010011000000000010100010000000000011010011000000000000000000000000000000000000000000");
		constant a_3 :std_logic_vector(107 downto 0) :=( "000000000000000000000000011010011000000000010100010000000000011010011000000000000000000000000000000000000000");
		constant a_4 :std_logic_vector(107 downto 0) :=( "000000000000000000000011010011000000000010100010000000000011010011000000000000000000000000000000000000000000");
		constant a_5 :std_logic_vector(107 downto 0) :=( "000000000000000000000000011010011000000000010100010000000000011010011000000000000000000000000000000000000000");
		constant a_6 :std_logic_vector(107 downto 0) :=( "000000000000000000000000000000000000000011010011000000000010100010000000000011010011000000000000000000000000");
		constant a_7 :std_logic_vector(107 downto 0) :=( "000000000000000000000000000000000000000000011010011000000000010100010000000000011010011000000000000000000000");
		constant b_0 :std_logic_vector(107 downto 0) :=( "000000000000000000000000000000000000000011010011000000000010100010000000000010001010000000000011010011000000");
		constant b_1 :std_logic_vector(107 downto 0) :=( "000000000000000000000000000000000000000000011010011000000000010100010000000000010001010000000000011010011000");
		constant b_2 :std_logic_vector(107 downto 0) :=( "000011010011000000000010001010000000000010100010000000000011010011000000000000000000000000000000000000000000");
		constant b_3 :std_logic_vector(107 downto 0) :=( "000000011010011000000000010001010000000000010100010000000000011010011000000000000000000000000000000000000000");
		constant b_4 :std_logic_vector(107 downto 0) :=( "000000000000000000011010010011000000010001100010000000011010010011000000000000000000000000000000000000000000");
		constant b_5 :std_logic_vector(107 downto 0) :=( "000000000000000000000000011010010011000000010100001010000000011010010011000000000000000000000000000000000000");
		constant b_6 :std_logic_vector(107 downto 0) :=( "000000000000000000000000000000000000011010010011000000010001100010000000011010010011000000000000000000000000");
		constant b_7 :std_logic_vector(107 downto 0) :=( "000000000000000000000000000000000000000000011010010011000000010100001010000000011010010011000000000000000000");
		constant c_0 :std_logic_vector(107 downto 0) :=( "000000000000000000000011010011000000000010001010000000000010100010000000000010001010000000000011010011000000");
		constant c_1 :std_logic_vector(107 downto 0) :=( "000000000000000000000000011010011000000000010001010000000000010100010000000000010001010000000000011010011000");
		constant c_2 :std_logic_vector(107 downto 0) :=( "000011010011000000000010001010000000000010100010000000000010001010000000000011010011000000000000000000000000");
		constant c_3 :std_logic_vector(107 downto 0) :=( "000000011010011000000000010001010000000000010100010000000000010001010000000000011010011000000000000000000000");
		constant c_4 :std_logic_vector(107 downto 0) :=( "000000000000000000011010010010011000010001100001010000011010010010011000000000000000000000000000000000000000");
		constant c_5 :std_logic_vector(107 downto 0) :=( "000000000000000000000011010010010011000010001100001010000011010010010011000000000000000000000000000000000000");
		constant c_6 :std_logic_vector(107 downto 0) :=( "000000000000000000000000000000000000011010010010011000010001100001010000011010010010011000000000000000000000");
		constant c_7 :std_logic_vector(107 downto 0) :=( "000000000000000000000000000000000000000011010010010011000010001100001010000011010010010011000000000000000000");
		constant d_0 :std_logic_vector(107 downto 0) :=( "000000000000000000000011010011000000000010001010011000000010100001010000000011010010011000000000000000000000");
		constant d_1 :std_logic_vector(107 downto 0) :=( "000000000000000000000000011010011000000011010001010000000010001100010000000011010010011000000000000000000000");
		constant d_2 :std_logic_vector(107 downto 0) :=( "000000000000000000000011010010011000000010100001010000000010001010011000000011010011000000000000000000000000");
		constant d_3 :std_logic_vector(107 downto 0) :=( "000000000000000000000011010010011000000010001100010000000011010001010000000000011010011000000000000000000000");
		constant d_4 :std_logic_vector(107 downto 0) :=( "000000000000000000000011010010011000000010100001010000000010001010011000000011010011000000000000000000000000");
		constant d_5 :std_logic_vector(107 downto 0) :=( "000000000000000000000011010010011000000010001100010000000011010001010000000000011010011000000000000000000000");
		constant d_6 :std_logic_vector(107 downto 0) :=( "000000000000000000000011010011000000000010001010011000000010100001010000000011010010011000000000000000000000");
		constant d_7 :std_logic_vector(107 downto 0) :=( "000000000000000000000000011010011000000011010001010000000010001100010000000011010010011000000000000000000000");
		constant e_0 :std_logic_vector(107 downto 0) :=( "000000000000000000000011010011000000000010001010000000011010100010000000010001001010000000011010010011000000");
		constant e_1 :std_logic_vector(107 downto 0) :=( "000000000000000000000000011010011000000000010001010000000000010100010011000000010001001010000000011010010011");
		constant e_2 :std_logic_vector(107 downto 0) :=( "011010010011000000010001001010000000011010100010000000000010001010000000000011010011000000000000000000000000");
		constant e_3 :std_logic_vector(107 downto 0) :=( "000000011010010011000000010001001010000000010100010011000000010001010000000000011010011000000000000000000000");
		constant e_4 :std_logic_vector(107 downto 0) :=( "011010011000000000010001010010011000010001100001010000011010010010011000000000000000000000000000000000000000");
		constant e_5 :std_logic_vector(107 downto 0) :=( "000000000011010011000011010010001010000010001100001010000011010010010011000000000000000000000000000000000000");
		constant e_6 :std_logic_vector(107 downto 0) :=( "000000000000000000000000000000000000011010010010011000010001100001010000010001010010011000011010011000000000");
		constant e_7 :std_logic_vector(107 downto 0) :=( "000000000000000000000000000000000000000011010010010011000010001100001010000011010010001010000000000011010011");
		constant f_0 :std_logic_vector(107 downto 0) :=( "000000000000000000000011010011000000000010001010011000000010100001010000000010001010011000000011010011000000");
		constant f_1 :std_logic_vector(107 downto 0) :=( "000000000000000000000000011010011000000011010001010000000010001100010000000011010001010000000000011010011000");
		constant f_2 :std_logic_vector(107 downto 0) :=( "000011010011000000000010001010011000000010100001010000000010001010011000000011010011000000000000000000000000");
		constant f_3 :std_logic_vector(107 downto 0) :=( "000000011010011000000011010001010000000010001100010000000011010001010000000000011010011000000000000000000000");
		constant f_4 :std_logic_vector(107 downto 0) :=( "000000000000000000011010010010011000010001100001010000011010001010011000000011010011000000000000000000000000");
		constant f_5 :std_logic_vector(107 downto 0) :=( "000000000000000000000011010010010011000010001100001010000011010001010011000000011010011000000000000000000000");
		constant f_6 :std_logic_vector(107 downto 0) :=( "000000000000000000000011010011000000011010001010011000010001100001010000011010010010011000000000000000000000");
		constant f_7 :std_logic_vector(107 downto 0) :=( "000000000000000000000000011010011000000011010001010011000010001100001010000011010010010011000000000000000000");
		constant g_0 :std_logic_vector(107 downto 0) :=( "000000000000000000000000000000000000000011010010011000000010100001010000000010001001010000000011010010011000");
		constant g_1 :std_logic_vector(107 downto 0) :=( "000000000000000000000000000000000000000011010010011000000010001100010000000010001001010000000011010010011000");
		constant g_2 :std_logic_vector(107 downto 0) :=( "000011010010011000000010001001010000000010100001010000000011010010011000000000000000000000000000000000000000");
		constant g_3 :std_logic_vector(107 downto 0) :=( "000011010010011000000010001001010000000010001100010000000011010010011000000000000000000000000000000000000000");
		constant g_4 :std_logic_vector(107 downto 0) :=( "000000000000000000011010010011000000010001100010000000010001001010000000011010010011000000000000000000000000");
		constant g_5 :std_logic_vector(107 downto 0) :=( "000000000000000000000000011010010011000000010100001010000000010001001010000000011010010011000000000000000000");
		constant g_6 :std_logic_vector(107 downto 0) :=( "000000000000000000011010010011000000010001001010000000010001100010000000011010010011000000000000000000000000");
		constant g_7 :std_logic_vector(107 downto 0) :=( "000000000000000000000000011010010011000000010001001010000000010100001010000000011010010011000000000000000000");
		constant h_0 :std_logic_vector(107 downto 0) :=( "000000000000000000000000000000000000011010010011000000010001100010011000011010001001010000000011010010011000");
		constant h_1 :std_logic_vector(107 downto 0) :=( "000000000000000000000000000000000000000000011010010011000011010100001010000010001001010011000011010010011000");
		constant h_2 :std_logic_vector(107 downto 0) :=( "000011010010011000011010001001010000010001100010011000011010010011000000000000000000000000000000000000000000");
		constant h_3 :std_logic_vector(107 downto 0) :=( "000011010010011000000010001001010011000011010100001010000000011010010011000000000000000000000000000000000000");
		constant h_4 :std_logic_vector(107 downto 0) :=( "000011010011000000011010001010000000010001100010000000010001010011000000011010011000000000000000000000000000");
		constant h_5 :std_logic_vector(107 downto 0) :=( "000000011010011000000000010001010011000000010100001010000000011010001010000000000011010011000000000000000000");
		constant h_6 :std_logic_vector(107 downto 0) :=( "000000000000000000011010011000000000010001010011000000010001100010000000011010001010000000000011010011000000");
		constant h_7 :std_logic_vector(107 downto 0) :=( "000000000000000000000000000011010011000000011010001010000000010100001010000000010001010011000000011010011000");
		constant i_0 :std_logic_vector(107 downto 0) :=( "000011010011000000000010001010000000011010001010000000010001100010000000010001010011000000011010011000000000");
		constant i_1 :std_logic_vector(107 downto 0) :=( "000000011010011000000000010001010000000000010001010011000000010100001010000000011010001010000000000011010011");
		constant i_2 :std_logic_vector(107 downto 0) :=( "011010011000000000010001010011000000010001100010000000011010001010000000000010001010000000000011010011000000");
		constant i_3 :std_logic_vector(107 downto 0) :=( "000000000011010011000000011010001010000000010100001010000000010001010011000000010001010000000000011010011000");
		constant i_4 :std_logic_vector(107 downto 0) :=( "011010010011000000010001001010010011011010100001001010000011010010010011000000000000000000000000000000000000");
		constant i_5 :std_logic_vector(107 downto 0) :=( "000000011010010011011010010001001010010001001100010011011010010010011000000000000000000000000000000000000000");
		constant i_6 :std_logic_vector(107 downto 0) :=( "000000000000000000000000000000000000000011010010010011011010100001001010010001001010010011011010010011000000");
		constant i_7 :std_logic_vector(107 downto 0) :=( "000000000000000000000000000000000000011010010010011000010001001100010011011010010001001010000000011010010011");
		constant j_0 :std_logic_vector(107 downto 0) :=( "000000000000000000000011010011000000011010001010000000010001100010000000010001001010000000011010010011000000");
		constant j_1 :std_logic_vector(107 downto 0) :=( "000000000000000000000000011010011000000000010001010011000000010100001010000000010001001010000000011010010011");
		constant j_2 :std_logic_vector(107 downto 0) :=( "011010010011000000010001001010000000010001100010000000011010001010000000000011010011000000000000000000000000");
		constant j_3 :std_logic_vector(107 downto 0) :=( "000000011010010011000000010001001010000000010100001010000000010001010011000000011010011000000000000000000000");
		constant j_4 :std_logic_vector(107 downto 0) :=( "011010010011000000010001001010011000010001100001010000011010010010011000000000000000000000000000000000000000");
		constant j_5 :std_logic_vector(107 downto 0) :=( "000000011010010011000011010001001010000010001100001010000011010010010011000000000000000000000000000000000000");
		constant j_6 :std_logic_vector(107 downto 0) :=( "000000000000000000000000000000000000011010010010011000010001100001010000010001001010011000011010010011000000");
		constant j_7 :std_logic_vector(107 downto 0) :=( "000000000000000000000000000000000000000011010010010011000010001100001010000011010001001010000000011010010011");
		constant k_0 :std_logic_vector(107 downto 0) :=( "000000000000000000011010010011000000010001001010000000011010100010000000010001001010000000011010010011000000");
		constant k_1 :std_logic_vector(107 downto 0) :=( "000000000000000000000000011010010011000000010001001010000000010100010011000000010001001010000000011010010011");
		constant k_2 :std_logic_vector(107 downto 0) :=( "011010010011000000010001001010000000011010100010000000010001001010000000011010010011000000000000000000000000");
		constant k_3 :std_logic_vector(107 downto 0) :=( "000000011010010011000000010001001010000000010100010011000000010001001010000000011010010011000000000000000000");
		constant k_4 :std_logic_vector(107 downto 0) :=( "011010011010011000010001010001010000010001100001010000011010010010011000000000000000000000000000000000000000");
		constant k_5 :std_logic_vector(107 downto 0) :=( "000011010011010011000010001010001010000010001100001010000011010010010011000000000000000000000000000000000000");
		constant k_6 :std_logic_vector(107 downto 0) :=( "000000000000000000000000000000000000011010010010011000010001100001010000010001010001010000011010011010011000");
		constant k_7 :std_logic_vector(107 downto 0) :=( "000000000000000000000000000000000000000011010010010011000010001100001010000010001010001010000011010011010011");
		constant l_0 :std_logic_vector(107 downto 0) :=( "000000000000000000000011010011000000000010001010000000011010100010011000010001001001010000011010010010011000");
		constant l_1 :std_logic_vector(107 downto 0) :=( "000000000000000000000000011010011000000000010001010000000011010100010011000010001001001010000011010010010011");
		constant l_2 :std_logic_vector(107 downto 0) :=( "011010010010011000010001001001010000011010100010011000000010001010000000000011010011000000000000000000000000");
		constant l_3 :std_logic_vector(107 downto 0) :=( "000011010010010011000010001001001010000011010100010011000000010001010000000000011010011000000000000000000000");
		constant l_4 :std_logic_vector(107 downto 0) :=( "011010011000000000010001010010011000010001100001010000010001010010011000011010011000000000000000000000000000");
		constant l_5 :std_logic_vector(107 downto 0) :=( "000000000011010011000011010010001010000010001100001010000011010010001010000000000011010011000000000000000000");
		constant l_6 :std_logic_vector(107 downto 0) :=( "000000000000000000011010011000000000010001010010011000010001100001010000010001010010011000011010011000000000");
		constant l_7 :std_logic_vector(107 downto 0) :=( "000000000000000000000000000011010011000011010010001010000010001100001010000011010010001010000000000011010011");
		constant m_0 :std_logic_vector(107 downto 0) :=( "000011010011000000000010001010000000000010001010010011000010100001001010000011010010010011000000000000000000");
		constant m_1 :std_logic_vector(107 downto 0) :=( "000000011010011000000000010001010000011010010001010000010001001100010000011010010010011000000000000000000000");
		constant m_2 :std_logic_vector(107 downto 0) :=( "000000000000000000000011010010010011000010100001001010000010001010010011000010001010000000000011010011000000");
		constant m_3 :std_logic_vector(107 downto 0) :=( "000000000000000000011010010010011000010001001100010000011010010001010000000000010001010000000000011010011000");
		constant m_4 :std_logic_vector(107 downto 0) :=( "000000000000000000000011010010010011000010100001001010000010001010010011000010001010000000000011010011000000");
		constant m_5 :std_logic_vector(107 downto 0) :=( "000000000000000000011010010010011000010001001100010000011010010001010000000000010001010000000000011010011000");
		constant m_6 :std_logic_vector(107 downto 0) :=( "000011010011000000000010001010000000000010001010010011000010100001001010000011010010010011000000000000000000");
		constant m_7 :std_logic_vector(107 downto 0) :=( "000000011010011000000000010001010000011010010001010000010001001100010000011010010010011000000000000000000000");
		constant n_0 :std_logic_vector(107 downto 0) :=( "000000000000000000011010010011000000010001001010011000011010100001010000000011010001010000000000011010011000");
		constant n_1 :std_logic_vector(107 downto 0) :=( "000000000000000000000000011010010011000011010001001010000010001100010011000010001010011000000011010011000000");
		constant n_2 :std_logic_vector(107 downto 0) :=( "000000011010011000000011010001010000011010100001010000010001001010011000011010010011000000000000000000000000");
		constant n_3 :std_logic_vector(107 downto 0) :=( "000011010011000000000010001010011000000010001100010011000011010001001010000000011010010011000000000000000000");
		constant n_4 :std_logic_vector(107 downto 0) :=( "000000011010011000000011010001010000011010100001010000010001001010011000011010010011000000000000000000000000");
		constant n_5 :std_logic_vector(107 downto 0) :=( "000011010011000000000010001010011000000010001100010011000011010001001010000000011010010011000000000000000000");
		constant n_6 :std_logic_vector(107 downto 0) :=( "000000000000000000011010010011000000010001001010011000011010100001010000000011010001010000000000011010011000");
		constant n_7 :std_logic_vector(107 downto 0) :=( "000000000000000000000000011010010011000011010001001010000010001100010011000010001010011000000011010011000000");
		constant o_0 :std_logic_vector(107 downto 0) :=( "000000000000000000011010011000000000010001010010011000010001100001010000011010010001010000000000011010011000");
		constant o_1 :std_logic_vector(107 downto 0) :=( "000000000000000000000000000011010011000011010010001010000010001100001010000010001010010011000011010011000000");
		constant o_2 :std_logic_vector(107 downto 0) :=( "000000011010011000011010010001010000010001100001010000010001010010011000011010011000000000000000000000000000");
		constant o_3 :std_logic_vector(107 downto 0) :=( "000011010011000000000010001010010011000010001100001010000011010010001010000000000011010011000000000000000000");
		constant o_4 :std_logic_vector(107 downto 0) :=( "000011010010011000000010001001010000011010100010011000010001001010000000011010010011000000000000000000000000");
		constant o_5 :std_logic_vector(107 downto 0) :=( "000011010010011000000010001001010000000011010100010011000000010001001010000000011010010011000000000000000000");
		constant o_6 :std_logic_vector(107 downto 0) :=( "000000000000000000011010010011000000010001001010000000011010100010011000000010001001010000000011010010011000");
		constant o_7 :std_logic_vector(107 downto 0) :=( "000000000000000000000000011010010011000000010001001010000011010100010011000010001001010000000011010010011000");
		constant p_0 :std_logic_vector(107 downto 0) :=( "000000000000000000011010011000000000010001010010011000010001100001010000011010001010011000000011010011000000");
		constant p_1 :std_logic_vector(107 downto 0) :=( "000000000000000000000000000011010011000011010010001010000010001100001010000011010001010011000000011010011000");
		constant p_2 :std_logic_vector(107 downto 0) :=( "000011010011000000011010001010011000010001100001010000010001010010011000011010011000000000000000000000000000");
		constant p_3 :std_logic_vector(107 downto 0) :=( "000000011010011000000011010001010011000010001100001010000011010010001010000000000011010011000000000000000000");
		constant p_4 :std_logic_vector(107 downto 0) :=( "000011010010011000011010001001010000010001100010011000011010001010000000000011010011000000000000000000000000");
		constant p_5 :std_logic_vector(107 downto 0) :=( "000011010010011000000010001001010011000011010100001010000000010001010011000000011010011000000000000000000000");
		constant p_6 :std_logic_vector(107 downto 0) :=( "000000000000000000000011010011000000011010001010000000010001100010011000011010001001010000000011010010011000");
		constant p_7 :std_logic_vector(107 downto 0) :=( "000000000000000000000000011010011000000000010001010011000011010100001010000010001001010011000011010010011000");
		constant q_0 :std_logic_vector(107 downto 0) :=( "000000000000000000000011010011000000011010001010011000010001100001010000011010001010011000000011010011000000");
		constant q_1 :std_logic_vector(107 downto 0) :=( "000000000000000000000000011010011000000011010001010011000010001100001010000011010001010011000000011010011000");
		constant q_2 :std_logic_vector(107 downto 0) :=( "000011010011000000011010001010011000010001100001010000011010001010011000000011010011000000000000000000000000");
		constant q_3 :std_logic_vector(107 downto 0) :=( "000000011010011000000011010001010011000010001100001010000011010001010011000000011010011000000000000000000000");
		constant q_4 :std_logic_vector(107 downto 0) :=( "000011010011000000011010001010011000010001100001010000011010001010011000000011010011000000000000000000000000");
		constant q_5 :std_logic_vector(107 downto 0) :=( "000000011010011000000011010001010011000010001100001010000011010001010011000000011010011000000000000000000000");
		constant q_6 :std_logic_vector(107 downto 0) :=( "000000000000000000000011010011000000011010001010011000010001100001010000011010001010011000000011010011000000");
		constant q_7 :std_logic_vector(107 downto 0) :=(	"000000000000000000000000011010011000000011010001010011000010001100001010000011010001010011000000011010011000");




begin



		sampler <= datain(107 downto 0);



--		 a(0)  <= ( "000000000000000000"&"000000000000000000"&"000011010011000000"&"000010100010000000"&"000011010011000000"&"000000000000000000");
--		 a(1)  <= (	"000000000000000000"&"000000000000000000"&"000000011010011000"&"000000010100010000"&"000000011010011000"&"000000000000000000");
--		 a(2)  <= ( "000000000000000000"&"000011010011000000"&"000010100010000000"&"000011010011000000"&"000000000000000000"&"000000000000000000");
--		 a(3)  <= ( "000000000000000000"&"000000011010011000"&"000000010100010000"&"000000011010011000"&"000000000000000000"&"000000000000000000");
--		 a(4)  <= ( "000000000000000000"&"000011010011000000"&"000010100010000000"&"000011010011000000"&"000000000000000000"&"000000000000000000");
--		 a(5)  <= ( "000000000000000000"&"000000011010011000"&"000000010100010000"&"000000011010011000"&"000000000000000000"&"000000000000000000");
--		 a(6)  <= ( "000000000000000000"&"000000000000000000"&"000011010011000000"&"000010100010000000"&"000011010011000000"&"000000000000000000");
--		 a(7)  <= ( "000000000000000000"&"000000000000000000"&"000000011010011000"&"000000010100010000"&"000000011010011000"&"000000000000000000");
--		 b(0)  <= ( "000000000000000000"&"000000000000000000"&"000011010011000000"&"000010100010000000"&"000010001010000000"&"000011010011000000");
--		 b(1)  <= ( "000000000000000000"&"000000000000000000"&"000000011010011000"&"000000010100010000"&"000000010001010000"&"000000011010011000");
--		 b(2)  <= ( "000011010011000000"&"000010001010000000"&"000010100010000000"&"000011010011000000"&"000000000000000000"&"000000000000000000");
--		 b(3)  <= ( "000000011010011000"&"000000010001010000"&"000000010100010000"&"000000011010011000"&"000000000000000000"&"000000000000000000");
--		 b(4)  <= ( "000000000000000000"&"011010010011000000"&"010001100010000000"&"011010010011000000"&"000000000000000000"&"000000000000000000");
--		 b(5)  <= ( "000000000000000000"&"000000011010010011"&"000000010100001010"&"000000011010010011"&"000000000000000000"&"000000000000000000");
--		 b(6)  <= ( "000000000000000000"&"000000000000000000"&"011010010011000000"&"010001100010000000"&"011010010011000000"&"000000000000000000");
--		 b(7)  <= ( "000000000000000000"&"000000000000000000"&"000000011010010011"&"000000010100001010"&"000000011010010011"&"000000000000000000");
--		 c(0)  <= ( "000000000000000000"&"000011010011000000"&"000010001010000000"&"000010100010000000"&"000010001010000000"&"000011010011000000");
--		 c(1)  <= ( "000000000000000000"&"000000011010011000"&"000000010001010000"&"000000010100010000"&"000000010001010000"&"000000011010011000");
--		 c(2)  <= ( "000011010011000000"&"000010001010000000"&"000010100010000000"&"000010001010000000"&"000011010011000000"&"000000000000000000");
--		 c(3)  <= ( "000000011010011000"&"000000010001010000"&"000000010100010000"&"000000010001010000"&"000000011010011000"&"000000000000000000");
--		 c(4)  <= ( "000000000000000000"&"011010010010011000"&"010001100001010000"&"011010010010011000"&"000000000000000000"&"000000000000000000");
--		 c(5)  <= ( "000000000000000000"&"000011010010010011"&"000010001100001010"&"000011010010010011"&"000000000000000000"&"000000000000000000");
--		 c(6)  <= ( "000000000000000000"&"000000000000000000"&"011010010010011000"&"010001100001010000"&"011010010010011000"&"000000000000000000");
--		 c(7)  <= ( "000000000000000000"&"000000000000000000"&"000011010010010011"&"000010001100001010"&"000011010010010011"&"000000000000000000");
--		 d(0)  <= ( "000000000000000000"&"000011010011000000"&"000010001010011000"&"000010100001010000"&"000011010010011000"&"000000000000000000");
--		 d(1)  <= ( "000000000000000000"&"000000011010011000"&"000011010001010000"&"000010001100010000"&"000011010010011000"&"000000000000000000");
--		 d(2)  <= ( "000000000000000000"&"000011010010011000"&"000010100001010000"&"000010001010011000"&"000011010011000000"&"000000000000000000");
--		 d(3)  <= ( "000000000000000000"&"000011010010011000"&"000010001100010000"&"000011010001010000"&"000000011010011000"&"000000000000000000");
--		 d(4)  <= ( "000000000000000000"&"000011010010011000"&"000010100001010000"&"000010001010011000"&"000011010011000000"&"000000000000000000");
--		 d(5)  <= ( "000000000000000000"&"000011010010011000"&"000010001100010000"&"000011010001010000"&"000000011010011000"&"000000000000000000");
--		 d(6)  <= ( "000000000000000000"&"000011010011000000"&"000010001010011000"&"000010100001010000"&"000011010010011000"&"000000000000000000");
--		 d(7)  <= ( "000000000000000000"&"000000011010011000"&"000011010001010000"&"000010001100010000"&"000011010010011000"&"000000000000000000");
--		 e(0)  <= ( "000000000000000000"&"000011010011000000"&"000010001010000000"&"011010100010000000"&"010001001010000000"&"011010010011000000");
--		 e(1)  <= ( "000000000000000000"&"000000011010011000"&"000000010001010000"&"000000010100010011"&"000000010001001010"&"000000011010010011");
--		 e(2)  <= ( "011010010011000000"&"010001001010000000"&"011010100010000000"&"000010001010000000"&"000011010011000000"&"000000000000000000");
--		 e(3)  <= ( "000000011010010011"&"000000010001001010"&"000000010100010011"&"000000010001010000"&"000000011010011000"&"000000000000000000");
--		 e(4)  <= ( "011010011000000000"&"010001010010011000"&"010001100001010000"&"011010010010011000"&"000000000000000000"&"000000000000000000");
--		 e(5)  <= ( "000000000011010011"&"000011010010001010"&"000010001100001010"&"000011010010010011"&"000000000000000000"&"000000000000000000");
--		 e(6)  <= ( "000000000000000000"&"000000000000000000"&"011010010010011000"&"010001100001010000"&"010001010010011000"&"011010011000000000");
--		 e(7)  <= ( "000000000000000000"&"000000000000000000"&"000011010010010011"&"000010001100001010"&"000011010010001010"&"000000000011010011");
--		 f(0)  <= ( "000000000000000000"&"000011010011000000"&"000010001010011000"&"000010100001010000"&"000010001010011000"&"000011010011000000");
--		 f(1)  <= ( "000000000000000000"&"000000011010011000"&"000011010001010000"&"000010001100010000"&"000011010001010000"&"000000011010011000");
--		 f(2)  <= ( "000011010011000000"&"000010001010011000"&"000010100001010000"&"000010001010011000"&"000011010011000000"&"000000000000000000");
--		 f(3)  <= ( "000000011010011000"&"000011010001010000"&"000010001100010000"&"000011010001010000"&"000000011010011000"&"000000000000000000");
--		 f(4)  <= ( "000000000000000000"&"011010010010011000"&"010001100001010000"&"011010001010011000"&"000011010011000000"&"000000000000000000");
--		 f(5)  <= ( "000000000000000000"&"000011010010010011"&"000010001100001010"&"000011010001010011"&"000000011010011000"&"000000000000000000");
--		 f(6)  <= ( "000000000000000000"&"000011010011000000"&"011010001010011000"&"010001100001010000"&"011010010010011000"&"000000000000000000");
--		 f(7)  <= ( "000000000000000000"&"000000011010011000"&"000011010001010011"&"000010001100001010"&"000011010010010011"&"000000000000000000");
--		 g(0)  <= ( "000000000000000000"&"000000000000000000"&"000011010010011000"&"000010100001010000"&"000010001001010000"&"000011010010011000");
--		 g(1)  <= ( "000000000000000000"&"000000000000000000"&"000011010010011000"&"000010001100010000"&"000010001001010000"&"000011010010011000");
--		 g(2)  <= ( "000011010010011000"&"000010001001010000"&"000010100001010000"&"000011010010011000"&"000000000000000000"&"000000000000000000");
--		 g(3)  <= ( "000011010010011000"&"000010001001010000"&"000010001100010000"&"000011010010011000"&"000000000000000000"&"000000000000000000");
--		 g(4)  <= ( "000000000000000000"&"011010010011000000"&"010001100010000000"&"010001001010000000"&"011010010011000000"&"000000000000000000");
--		 g(5)  <= ( "000000000000000000"&"000000011010010011"&"000000010100001010"&"000000010001001010"&"000000011010010011"&"000000000000000000");
--		 g(6)  <= ( "000000000000000000"&"011010010011000000"&"010001001010000000"&"010001100010000000"&"011010010011000000"&"000000000000000000");
--		 g(7)  <= ( "000000000000000000"&"000000011010010011"&"000000010001001010"&"000000010100001010"&"000000011010010011"&"000000000000000000");
--		 h(0)  <= ( "000000000000000000"&"000000000000000000"&"011010010011000000"&"010001100010011000"&"011010001001010000"&"000011010010011000");
--		 h(1)  <= ( "000000000000000000"&"000000000000000000"&"000000011010010011"&"000011010100001010"&"000010001001010011"&"000011010010011000");
--		 h(2)  <= ( "000011010010011000"&"011010001001010000"&"010001100010011000"&"011010010011000000"&"000000000000000000"&"000000000000000000");
--		 h(3)  <= ( "000011010010011000"&"000010001001010011"&"000011010100001010"&"000000011010010011"&"000000000000000000"&"000000000000000000");
--		 h(4)  <= ( "000011010011000000"&"011010001010000000"&"010001100010000000"&"010001010011000000"&"011010011000000000"&"000000000000000000");
--		 h(5)  <= ( "000000011010011000"&"000000010001010011"&"000000010100001010"&"000000011010001010"&"000000000011010011"&"000000000000000000");
--		 h(6)  <= ( "000000000000000000"&"011010011000000000"&"010001010011000000"&"010001100010000000"&"011010001010000000"&"000011010011000000");
--		 h(7)  <= ( "000000000000000000"&"000000000011010011"&"000000011010001010"&"000000010100001010"&"000000010001010011"&"000000011010011000");
--		 i(0)  <= ( "000011010011000000"&"000010001010000000"&"011010001010000000"&"010001100010000000"&"010001010011000000"&"011010011000000000");
--		 i(1)  <= ( "000000011010011000"&"000000010001010000"&"000000010001010011"&"000000010100001010"&"000000011010001010"&"000000000011010011");
--		 i(2)  <= ( "011010011000000000"&"010001010011000000"&"010001100010000000"&"011010001010000000"&"000010001010000000"&"000011010011000000");
--		 i(3)  <= ( "000000000011010011"&"000000011010001010"&"000000010100001010"&"000000010001010011"&"000000010001010000"&"000000011010011000");
--		 i(4)  <= ( "011010010011000000"&"010001001010010011"&"011010100001001010"&"000011010010010011"&"000000000000000000"&"000000000000000000");
--		 i(5)  <= ( "000000011010010011"&"011010010001001010"&"010001001100010011"&"011010010010011000"&"000000000000000000"&"000000000000000000");
--		 i(6)  <= ( "000000000000000000"&"000000000000000000"&"000011010010010011"&"011010100001001010"&"010001001010010011"&"011010010011000000");
--		 i(7)  <= ( "000000000000000000"&"000000000000000000"&"011010010010011000"&"010001001100010011"&"011010010001001010"&"000000011010010011");
--		 j(0)  <= ( "000000000000000000"&"000011010011000000"&"011010001010000000"&"010001100010000000"&"010001001010000000"&"011010010011000000");
--		 j(1)  <= ( "000000000000000000"&"000000011010011000"&"000000010001010011"&"000000010100001010"&"000000010001001010"&"000000011010010011");
--		 j(2)  <= ( "011010010011000000"&"010001001010000000"&"010001100010000000"&"011010001010000000"&"000011010011000000"&"000000000000000000");
--		 j(3)  <= ( "000000011010010011"&"000000010001001010"&"000000010100001010"&"000000010001010011"&"000000011010011000"&"000000000000000000");
--		 j(4)  <= ( "011010010011000000"&"010001001010011000"&"010001100001010000"&"011010010010011000"&"000000000000000000"&"000000000000000000");
--		 j(5)  <= ( "000000011010010011"&"000011010001001010"&"000010001100001010"&"000011010010010011"&"000000000000000000"&"000000000000000000");
--		 j(6)  <= ( "000000000000000000"&"000000000000000000"&"011010010010011000"&"010001100001010000"&"010001001010011000"&"011010010011000000");
--		 j(7)  <= ( "000000000000000000"&"000000000000000000"&"000011010010010011"&"000010001100001010"&"000011010001001010"&"000000011010010011");
--		 k(0)  <= ( "000000000000000000"&"011010010011000000"&"010001001010000000"&"011010100010000000"&"010001001010000000"&"011010010011000000");
--		 k(1)  <= ( "000000000000000000"&"000000011010010011"&"000000010001001010"&"000000010100010011"&"000000010001001010"&"000000011010010011");
--		 k(2)  <= ( "011010010011000000"&"010001001010000000"&"011010100010000000"&"010001001010000000"&"011010010011000000"&"000000000000000000");
--		 k(3)  <= ( "000000011010010011"&"000000010001001010"&"000000010100010011"&"000000010001001010"&"000000011010010011"&"000000000000000000");
--		 k(4)  <= ( "011010011010011000"&"010001010001010000"&"010001100001010000"&"011010010010011000"&"000000000000000000"&"000000000000000000");
--		 k(5)  <= ( "000011010011010011"&"000010001010001010"&"000010001100001010"&"000011010010010011"&"000000000000000000"&"000000000000000000");
--		 k(6)  <= ( "000000000000000000"&"000000000000000000"&"011010010010011000"&"010001100001010000"&"010001010001010000"&"011010011010011000");
--		 k(7)  <= ( "000000000000000000"&"000000000000000000"&"000011010010010011"&"000010001100001010"&"000010001010001010"&"000011010011010011");
--		 l(0)  <= ( "000000000000000000"&"000011010011000000"&"000010001010000000"&"011010100010011000"&"010001001001010000"&"011010010010011000");
--		 l(1)  <= ( "000000000000000000"&"000000011010011000"&"000000010001010000"&"000011010100010011"&"000010001001001010"&"000011010010010011");
--		 l(2)  <= ( "011010010010011000"&"010001001001010000"&"011010100010011000"&"000010001010000000"&"000011010011000000"&"000000000000000000");
--		 l(3)  <= ( "000011010010010011"&"000010001001001010"&"000011010100010011"&"000000010001010000"&"000000011010011000"&"000000000000000000");
--		 l(4)  <= ( "011010011000000000"&"010001010010011000"&"010001100001010000"&"010001010010011000"&"011010011000000000"&"000000000000000000");
--		 l(5)  <= ( "000000000011010011"&"000011010010001010"&"000010001100001010"&"000011010010001010"&"000000000011010011"&"000000000000000000");
--		 l(6)  <= ( "000000000000000000"&"011010011000000000"&"010001010010011000"&"010001100001010000"&"010001010010011000"&"011010011000000000");
--		 l(7)  <= ( "000000000000000000"&"000000000011010011"&"000011010010001010"&"000010001100001010"&"000011010010001010"&"000000000011010011");
--		 m(0)  <= ( "000011010011000000"&"000010001010000000"&"000010001010010011"&"000010100001001010"&"000011010010010011"&"000000000000000000");
--		 m(1)  <= ( "000000011010011000"&"000000010001010000"&"011010010001010000"&"010001001100010000"&"011010010010011000"&"000000000000000000");
--		 m(2)  <= ( "000000000000000000"&"000011010010010011"&"000010100001001010"&"000010001010010011"&"000010001010000000"&"000011010011000000");
--		 m(3)  <= ( "000000000000000000"&"011010010010011000"&"010001001100010000"&"011010010001010000"&"000000010001010000"&"000000011010011000");
--		 m(4)  <= ( "000000000000000000"&"000011010010010011"&"000010100001001010"&"000010001010010011"&"000010001010000000"&"000011010011000000");
--		 m(5)  <= ( "000000000000000000"&"011010010010011000"&"010001001100010000"&"011010010001010000"&"000000010001010000"&"000000011010011000");
--		 m(6)  <= ( "000011010011000000"&"000010001010000000"&"000010001010010011"&"000010100001001010"&"000011010010010011"&"000000000000000000");
--		 m(7)  <= ( "000000011010011000"&"000000010001010000"&"011010010001010000"&"010001001100010000"&"011010010010011000"&"000000000000000000");
--		 n(0)  <= ( "000000000000000000"&"011010010011000000"&"010001001010011000"&"011010100001010000"&"000011010001010000"&"000000011010011000");
--		 n(1)  <= ( "000000000000000000"&"000000011010010011"&"000011010001001010"&"000010001100010011"&"000010001010011000"&"000011010011000000");
--		 n(2)  <= ( "000000011010011000"&"000011010001010000"&"011010100001010000"&"010001001010011000"&"011010010011000000"&"000000000000000000");
--		 n(3)  <= ( "000011010011000000"&"000010001010011000"&"000010001100010011"&"000011010001001010"&"000000011010010011"&"000000000000000000");
--		 n(4)  <= ( "000000011010011000"&"000011010001010000"&"011010100001010000"&"010001001010011000"&"011010010011000000"&"000000000000000000");
--		 n(5)  <= ( "000011010011000000"&"000010001010011000"&"000010001100010011"&"000011010001001010"&"000000011010010011"&"000000000000000000");
--		 n(6)  <= ( "000000000000000000"&"011010010011000000"&"010001001010011000"&"011010100001010000"&"000011010001010000"&"000000011010011000");
--		 n(7)  <= ( "000000000000000000"&"000000011010010011"&"000011010001001010"&"000010001100010011"&"000010001010011000"&"000011010011000000");
--		 o(0)  <= ( "000000000000000000"&"011010011000000000"&"010001010010011000"&"010001100001010000"&"011010010001010000"&"000000011010011000");
--		 o(1)  <= ( "000000000000000000"&"000000000011010011"&"000011010010001010"&"000010001100001010"&"000010001010010011"&"000011010011000000");
--		 o(2)  <= ( "000000011010011000"&"011010010001010000"&"010001100001010000"&"010001010010011000"&"011010011000000000"&"000000000000000000");
--		 o(3)  <= ( "000011010011000000"&"000010001010010011"&"000010001100001010"&"000011010010001010"&"000000000011010011"&"000000000000000000");
--		 o(4)  <= ( "000011010010011000"&"000010001001010000"&"011010100010011000"&"010001001010000000"&"011010010011000000"&"000000000000000000");
--		 o(5)  <= ( "000011010010011000"&"000010001001010000"&"000011010100010011"&"000000010001001010"&"000000011010010011"&"000000000000000000");
--		 o(6)  <= ( "000000000000000000"&"011010010011000000"&"010001001010000000"&"011010100010011000"&"000010001001010000"&"000011010010011000");
--		 o(7)  <= ( "000000000000000000"&"000000011010010011"&"000000010001001010"&"000011010100010011"&"000010001001010000"&"000011010010011000");
--		 p(0)  <= ( "000000000000000000"&"011010011000000000"&"010001010010011000"&"010001100001010000"&"011010001010011000"&"000011010011000000");
--		 p(1)  <= ( "000000000000000000"&"000000000011010011"&"000011010010001010"&"000010001100001010"&"000011010001010011"&"000000011010011000");
--		 p(2)  <= ( "000011010011000000"&"011010001010011000"&"010001100001010000"&"010001010010011000"&"011010011000000000"&"000000000000000000");
--		 p(3)  <= ( "000000011010011000"&"000011010001010011"&"000010001100001010"&"000011010010001010"&"000000000011010011"&"000000000000000000");
--		 p(4)  <= ( "000011010010011000"&"011010001001010000"&"010001100010011000"&"011010001010000000"&"000011010011000000"&"000000000000000000");
--		 p(5)  <= ( "000011010010011000"&"000010001001010011"&"000011010100001010"&"000000010001010011"&"000000011010011000"&"000000000000000000");
--		 p(6)  <= ( "000000000000000000"&"000011010011000000"&"011010001010000000"&"010001100010011000"&"011010001001010000"&"000011010010011000");
--		 p(7)  <= ( "000000000000000000"&"000000011010011000"&"000000010001010011"&"000011010100001010"&"000010001001010011"&"000011010010011000");
--		 q(0)  <= ( "000000000000000000"&"000011010011000000"&"011010001010011000"&"010001100001010000"&"011010001010011000"&"000011010011000000");
--		 q(1)  <= ( "000000000000000000"&"000000011010011000"&"000011010001010011"&"000010001100001010"&"000011010001010011"&"000000011010011000");
--		 q(2)  <= ( "000011010011000000"&"011010001010011000"&"010001100001010000"&"011010001010011000"&"000011010011000000"&"000000000000000000");
--		 q(3)  <= ( "000000011010011000"&"000011010001010011"&"000010001100001010"&"000011010001010011"&"000000011010011000"&"000000000000000000");
--		 q(4)  <= ( "000011010011000000"&"011010001010011000"&"010001100001010000"&"011010001010011000"&"000011010011000000"&"000000000000000000");
--		 q(5)  <= ( "000000011010011000"&"000011010001010011"&"000010001100001010"&"000011010001010011"&"000000011010011000"&"000000000000000000");
--		 q(6)  <= ( "000000000000000000"&"000011010011000000"&"011010001010011000"&"010001100001010000"&"011010001010011000"&"000011010011000000");
--		 q(7)  <= (	"000000000000000000"&"000000011010011000"&"000011010001010011"&"000010001100001010"&"000011010001010011"&"000000011010011000");


--		with sampler select
--			X_black_inner <= unsigned(datain(117 downto 113))- 3 when a(0)|a(2)|a(4)|a(6)|b(0)|b(2)|b(4)|b(6)|c(0)|c(2)|c(4)|c(6)|d(0)|d(2)|d(4)|d(6)|e(0)|e(2)|e(4)|e(6)|f(0)|f(2)|f(4)|f(6)|g(0)|g(2)|g(4)|g(6)|h(0)|h(2)|h(4)|h(6)|i(0)|i(2)|i(4)|i(6)|j(0)|j(2)|j(4)|j(6)|k(0)|k(2)|k(4)|k(6)|l(0)|l(2)|l(4)|l(6)|m(0)|m(2)|m(4)|m(6)|n(0)|n(2)|n(4)|n(6)|o(0)|o(2)|o(4)|o(6)|p(0)|p(2)|p(4)|p(6)|q(0)|q(2)|q(4)|q(6),
--								unsigned(datain(117 downto 113))- 2 when others;

		with sampler select
			X_black_before <= unsigned(datain(117 downto 113))- 3 when a_0|a_2|b_0|b_2|b_4|b_6|c_0|c_2|c_4|c_6|d_0|d_2|e_0|e_2|e_4|e_6|f_0|f_2|f_4|f_6|g_0|g_2|g_4|g_6|h_0|h_2|h_4|h_6|i_0|i_2|i_4|i_6|j_0|j_2|j_4|j_6|k_0|k_2|k_4|k_6|l_0|l_2|l_4|l_6|m_0|m_2|n_0|n_2|o_0|o_2|o_4|o_6|p_0|p_2|p_4|p_6|q_0|q_2,
								unsigned(datain(117 downto 113))- 2 when others;								

		--X_black_before <= 15 - X_black_inner;
--
--		with X_black_before select
--			X_black <= "01100011" when "01010",
--								"1100010" when "01011",
--								"1100011" when "01100",
--								("00" & X_black_before)  when others;						
--	
--
		with X_black_before select
			X_black <= "01100011" when "00011",
								"01100010" when "00100",
								"01100001" when "00101",
								"00111001" when "00110",
								"00111000" when	"00111",
								"00110111" when	"01000",
								"00110110" when	"01001",
								"00110101" when	"01010",
								"00110100" when	"01011",
								"00110011" when	"01100",
								"00110010" when	"01101",
								"00110001" when "01110",
								"00000000" when others;

--
--		with sampler select
--			Y_black_inner <= unsigned(datain(112 downto 108))-	2 when a(0)|a(1)|a(7)|a(6)|b(0)|b(1)|b(7)|b(6)|c(0)|c(1)|c(7)|c(6)|d(0)|d(1)|d(7)|d(6)|e(0)|e(1)|e(7)|e(6)|f(0)|f(1)|f(7)|f(6)|g(0)|g(1)|g(7)|g(6)|h(0)|h(1)|h(7)|h(6)|i(0)|i(1)|i(7)|i(6)|j(0)|j(1)|j(7)|j(6)|k(0)|k(1)|k(7)|k(6)|l(0)|l(1)|l(7)|l(6)|m(0)|m(1)|m(7)|m(6)|n(0)|n(1)|n(7)|n(6)|o(0)|o(1)|o(7)|o(6)|p(0)|p(1)|p(7)|p(6)|q(0)|q(1)|q(7)|q(6),
--								unsigned(datain(112 downto 108))-	3 when others;
--

		with sampler select
			Y_black_before <= unsigned(datain(112 downto 108))-	2 when a_0|a_1|b_0|b_1|b_7|b_6|c_0|c_1|c_7|c_6|d_0|d_1|e_0|e_1|e_7|e_6|f_0|f_1|f_7|f_6|g_0|g_1|g_7|g_6|h_0|h_1|h_7|h_6|i_0|i_1|i_7|i_6|j_0|j_1|j_7|j_6|k_0|k_1|k_7|k_6|l_0|l_1|l_7|l_6|m_0|m_1|n_0|n_1|o_0|o_1|o_7|o_6|p_0|p_1|p_7|p_6|q_0|q_1,
								unsigned(datain(112 downto 108))-	3 when others;


	--	Y_black_before <= 15 - Y_black_inner;
	--	Y_black_before <= "0001101";
		with Y_black_before select
			Y_black <= "01100011" when "00011",
								"01100010" when "00100",
								"01100001" when "00101",
								"00111001" when "00110",
								"00111000" when	"00111",
								"00110111" when	"01000",
								"00110110" when	"01001",
								"00110101" when	"01010",
								"00110100" when	"01011",
								"00110011" when	"01100",
								"00110010" when	"01101",
								"00110001" when "01110",
								"00000000" when others;

--		with sampler select
--			rotate <= "000" when a(0)|b(0)|c(0)|d(0)|e(0)|f(0)|g(0)|h(0)|i(0)|j(0)|k(0)|l(0)|m(0)|n(0)|o(0)|p(0)|q(0) ,
--								"001" when a(1)|b(1)|c(1)|d(1)|e(1)|f(1)|g(1)|h(1)|i(1)|j(1)|k(1)|l(1)|m(1)|n(1)|o(1)|p(1)|q(1) ,
--								"010" when a(2)|b(2)|c(2)|d(2)|e(2)|f(2)|g(2)|h(2)|i(2)|j(2)|k(2)|l(2)|m(2)|n(2)|o(2)|p(2)|q(2) ,
--								"011" when a(3)|b(3)|c(3)|d(3)|e(3)|f(3)|g(3)|h(3)|i(3)|j(3)|k(3)|l(3)|m(3)|n(3)|o(3)|p(3)|q(3) ,
--								"100" when a(4)|b(4)|c(4)|d(4)|e(4)|f(4)|g(4)|h(4)|i(4)|j(4)|k(4)|l(4)|m(4)|n(4)|o(4)|p(4)|q(4) ,
--								"101" when a(5)|b(5)|c(5)|d(5)|e(5)|f(5)|g(5)|h(5)|i(5)|j(5)|k(5)|l(5)|m(5)|n(5)|o(5)|p(5)|q(5) ,
--								"110" when a(6)|b(6)|c(6)|d(6)|e(6)|f(6)|g(6)|h(6)|i(6)|j(6)|k(6)|l(6)|m(6)|n(6)|o(6)|p(6)|q(6) ,
--								"111" when others;

		with sampler select
			rotate <= "00110000" when a_0|b_0|c_0|d_0|e_0|f_0|g_0|h_0|i_0|j_0|k_0|l_0|m_0|n_0|o_0|p_0|q_0 ,
								"00110001" when a_1|b_1|c_1|d_1|e_1|f_1|g_1|h_1|i_1|j_1|k_1|l_1|m_1|n_1|o_1|p_1|q_1 ,
								"00110010" when a_2|b_2|c_2|d_2|e_2|f_2|g_2|h_2|i_2|j_2|k_2|l_2|m_2|n_2|o_2|p_2|q_2 ,
								"00110011" when a_3|b_3|c_3|d_3|e_3|f_3|g_3|h_3|i_3|j_3|k_3|l_3|m_3|n_3|o_3|p_3|q_3 ,
								"00110100" when b_4|c_4|e_4|f_4|g_4|h_4|i_4|j_4|k_4|l_4|o_4|p_4 ,
								"00110101" when b_5|c_5|e_5|f_5|g_5|h_5|i_5|j_5|k_5|l_5|o_5|p_5 ,
								"00110110" when b_6|c_6|e_6|f_6|g_6|h_6|i_6|j_6|k_6|l_6|o_6|p_6 ,
								"00110111" when others;								
--
--		with sampler select
--			format <= "1100001" when a(0)|a(1)|a(2)|a(3)|a(4)|a(5)|a(6)|a(7) ,
--								"1100010" when b(0)|b(1)|b(2)|b(3)|b(4)|b(5)|b(6)|b(7) ,
--								"1100011" when c(0)|c(1)|c(2)|c(3)|c(4)|c(5)|c(6)|c(7) ,
--								"1100100" when d(0)|d(1)|d(2)|d(3)|d(4)|d(5)|d(6)|d(7) ,
--								"1100101" when e(0)|e(1)|e(2)|e(3)|e(4)|e(5)|e(6)|e(7) ,
--								"1100110" when f(0)|f(1)|f(2)|f(3)|f(4)|f(5)|f(6)|f(7) ,
--								"1100111" when g(0)|g(1)|g(2)|g(3)|g(4)|g(5)|g(6)|g(7) ,
--								"1101000" when h(0)|h(1)|h(2)|h(3)|h(4)|h(5)|h(6)|h(7) ,
--								"1101001" when i(0)|i(1)|i(2)|i(3)|i(4)|i(5)|i(6)|i(7) ,
--								"1101010" when j(0)|j(1)|j(2)|j(3)|j(4)|j(5)|j(6)|j(7) ,
--								"1101011" when k(0)|k(1)|k(2)|k(3)|k(4)|k(5)|k(6)|k(7) ,
--								"1101100" when l(0)|l(1)|l(2)|l(3)|l(4)|l(5)|l(6)|l(7) ,
--								"1101101" when m(0)|m(1)|m(2)|m(3)|m(4)|m(5)|m(6)|m(7) ,
--								"1101110" when n(0)|n(1)|n(2)|n(3)|n(4)|n(5)|n(6)|n(7) ,
--								"1101111" when o(0)|o(1)|o(2)|o(3)|o(4)|o(5)|o(6)|o(7),
--								"1110000" when p(0)|p(1)|p(2)|p(3)|p(4)|p(5)|p(6)|p(7) ,
--								"1110001" when others;

		with sampler select
			format <= "01100001" when a_0|a_1|a_2|a_3 ,
								"01100010" when b_0|b_1|b_2|b_3|b_4|b_5|b_6|b_7 ,
								"01100011" when c_0|c_1|c_2|c_3|c_4|c_5|c_6|c_7 ,
								"01100100" when d_0|d_1|d_2|d_3 ,
								"01100101" when e_0|e_1|e_2|e_3|e_4|e_5|e_6|e_7 ,
								"01100110" when f_0|f_1|f_2|f_3|f_4|f_5|f_6|f_7 ,
								"01100111" when g_0|g_1|g_2|g_3|g_4|g_5|g_6|g_7 ,
								"01101000" when h_0|h_1|h_2|h_3|h_4|h_5|h_6|h_7 ,
								"01101001" when i_0|i_1|i_2|i_3|i_4|i_5|i_6|i_7 ,
								"01101010" when j_0|j_1|j_2|j_3|j_4|j_5|j_6|j_7 ,
								"01101011" when k_0|k_1|k_2|k_3|k_4|k_5|k_6|k_7 ,
								"01101100" when l_0|l_1|l_2|l_3|l_4|l_5|l_6|l_7 ,
								"01101101" when m_0|m_1|m_2|m_3 ,
								"01101110" when n_0|n_1|n_2|n_3 ,
								"01101111" when o_0|o_1|o_2|o_3|o_4|o_5|o_6|o_7,
								"01110000" when p_0|p_1|p_2|p_3|p_4|p_5|p_6|p_7 ,
								"01110001" when others;
														

	data_coded <= (std_logic_vector(X_black) & std_logic_vector(Y_black) & std_logic_vector(format) & std_logic_vector(rotate));





end Gate_level;


---------------------------------------------------------------------------------------------------------------------------------
architecture test_bench of program_coding is

  -- Component Declaration
Component x Port (datain : in std_logic_vector (117 downto 0);
 								data_coded : out std_logic_vector(31 downto 0) 
				  );
end component;
for g:x use Entity work.program_coding(Gate_level);

signal datain1 : std_logic_vector(117 downto 0);
signal data_coded1 : std_logic_vector (31 downto 0);
begin

-- Component Instantiation
  g: x PORT MAP(datain1,data_coded1);
		 
    datain1 <= "0011101011000000000000000000000000000000000000000011010011000000000010100010000000000010001010000000000011010011000000"; --"1100000000000000" after 2 ns,"1010101010101010" after 4 ns,"1111111111111111" after 6 ns,"1111111100000000" after 8 ns,"1111110011001001" after 10 ns; '1','0' after 10 ns;

end test_bench;



