





library IEEE;
use IEEE.STD_logic_1164.ALL;
use IEEE.numeric_std.ALL;

entity  code is 
port (
data_code_ch : out std_logic;
load_code : in std_logic;
round : in std_logic_vector(1 downto 0);
data_rec : in std_logic;
ok : out std_logic_vector(117 downto 0);
load : out std_logic;
din : in std_logic_vector(117 downto 0);
clk : in std_logic);

end code;

architecture failure of code is 

type matrix is array (11 downto 0) of std_logic_vector(35 downto 0);
type  pieces is array (5 downto 0) of std_logic_vector(17 downto 0);
type generalmat is array (135 downto 0) of std_logic_vector(107 downto 0);
signal P,P_next,opp,opp_next: matrix := (others => (others => '0') );
signal aaa : matrix;
signal M,M_reg: pieces ;
-- signal state_reg,state_next : std_logic_vector(2 downto 0) := "000";
signal state_reg,state_next : std_logic_vector(1 downto 0);
--signal a: string (1 to 6) ;
signal sw1,sw2,sw1_next,sw2_next : std_logic := '0';
signal load_reg,load_next : std_logic := '0';	
signal form_next,form : std_logic_vector(15 downto 0) := (others => '0');	
signal formnex,formnex_next : std_logic_vector(15 downto 0) := (others => '0');	
signal rotate,rotate_next : std_logic_vector(7 downto 0) := (others => '0');
signal dout_reg , dout_next : std_logic_vector(117 downto 0);
signal x_reg,x_next,y_reg,y_next,x_in,y_in: integer range 0 to 20:= 0; -- for test bench 4
signal data_code_ch_reg,data_code_ch_next : std_logic := '0';

		constant a_0 :pieces :=( "000000000000000000","000000000000000000","000011010011000000","000010100010000000","000011010011000000","000000000000000000");
		constant a_1 :pieces :=(	"000000000000000000","000000000000000000","000000011010011000","000000010100010000","000000011010011000","000000000000000000");
		constant a_2 :pieces :=( "000000000000000000","000011010011000000","000010100010000000","000011010011000000","000000000000000000","000000000000000000");
		constant a_3 :pieces :=( "000000000000000000","000000011010011000","000000010100010000","000000011010011000","000000000000000000","000000000000000000");
		constant a_4 :pieces :=( "000000000000000000","000011010011000000","000010100010000000","000011010011000000","000000000000000000","000000000000000000");
		constant a_5 :pieces :=( "000000000000000000","000000011010011000","000000010100010000","000000011010011000","000000000000000000","000000000000000000");
		constant a_6 :pieces :=( "000000000000000000","000000000000000000","000011010011000000","000010100010000000","000011010011000000","000000000000000000");
		constant a_7 :pieces :=( "000000000000000000","000000000000000000","000000011010011000","000000010100010000","000000011010011000","000000000000000000");
		constant b_0 :pieces :=( "000000000000000000","000000000000000000","000011010011000000","000010100010000000","000010001010000000","000011010011000000");
		constant b_1 :pieces :=( "000000000000000000","000000000000000000","000000011010011000","000000010100010000","000000010001010000","000000011010011000");
		constant b_2 :pieces :=( "000011010011000000","000010001010000000","000010100010000000","000011010011000000","000000000000000000","000000000000000000");
		constant b_3 :pieces :=( "000000011010011000","000000010001010000","000000010100010000","000000011010011000","000000000000000000","000000000000000000");
		constant b_4 :pieces :=( "000000000000000000","011010010011000000","010001100010000000","011010010011000000","000000000000000000","000000000000000000");
		constant b_5 :pieces :=( "000000000000000000","000000011010010011","000000010100001010","000000011010010011","000000000000000000","000000000000000000");
		constant b_6 :pieces :=( "000000000000000000","000000000000000000","011010010011000000","010001100010000000","011010010011000000","000000000000000000");
		constant b_7 :pieces :=( "000000000000000000","000000000000000000","000000011010010011","000000010100001010","000000011010010011","000000000000000000");
		constant c_0 :pieces :=( "000000000000000000","000011010011000000","000010001010000000","000010100010000000","000010001010000000","000011010011000000");
		constant c_1 :pieces :=( "000000000000000000","000000011010011000","000000010001010000","000000010100010000","000000010001010000","000000011010011000");
		constant c_2 :pieces :=( "000011010011000000","000010001010000000","000010100010000000","000010001010000000","000011010011000000","000000000000000000");
		constant c_3 :pieces :=( "000000011010011000","000000010001010000","000000010100010000","000000010001010000","000000011010011000","000000000000000000");
		constant c_4 :pieces :=( "000000000000000000","011010010010011000","010001100001010000","011010010010011000","000000000000000000","000000000000000000");
		constant c_5 :pieces :=( "000000000000000000","000011010010010011","000010001100001010","000011010010010011","000000000000000000","000000000000000000");
		constant c_6 :pieces :=( "000000000000000000","000000000000000000","011010010010011000","010001100001010000","011010010010011000","000000000000000000");
		constant c_7 :pieces :=( "000000000000000000","000000000000000000","000011010010010011","000010001100001010","000011010010010011","000000000000000000");
		constant d_0 :pieces :=( "000000000000000000","000011010011000000","000010001010011000","000010100001010000","000011010010011000","000000000000000000");
		constant d_1 :pieces :=( "000000000000000000","000000011010011000","000011010001010000","000010001100010000","000011010010011000","000000000000000000");
		constant d_2 :pieces :=( "000000000000000000","000011010010011000","000010100001010000","000010001010011000","000011010011000000","000000000000000000");
		constant d_3 :pieces :=( "000000000000000000","000011010010011000","000010001100010000","000011010001010000","000000011010011000","000000000000000000");
		constant d_4 :pieces :=( "000000000000000000","000011010010011000","000010100001010000","000010001010011000","000011010011000000","000000000000000000");
		constant d_5 :pieces :=( "000000000000000000","000011010010011000","000010001100010000","000011010001010000","000000011010011000","000000000000000000");
		constant d_6 :pieces :=( "000000000000000000","000011010011000000","000010001010011000","000010100001010000","000011010010011000","000000000000000000");
		constant d_7 :pieces :=( "000000000000000000","000000011010011000","000011010001010000","000010001100010000","000011010010011000","000000000000000000");
		constant e_0 :pieces :=( "000000000000000000","000011010011000000","000010001010000000","011010100010000000","010001001010000000","011010010011000000");
		constant e_1 :pieces :=( "000000000000000000","000000011010011000","000000010001010000","000000010100010011","000000010001001010","000000011010010011");
		constant e_2 :pieces :=( "011010010011000000","010001001010000000","011010100010000000","000010001010000000","000011010011000000","000000000000000000");
		constant e_3 :pieces :=( "000000011010010011","000000010001001010","000000010100010011","000000010001010000","000000011010011000","000000000000000000");
		constant e_4 :pieces :=( "011010011000000000","010001010010011000","010001100001010000","011010010010011000","000000000000000000","000000000000000000");
		constant e_5 :pieces :=( "000000000011010011","000011010010001010","000010001100001010","000011010010010011","000000000000000000","000000000000000000");
		constant e_6 :pieces :=( "000000000000000000","000000000000000000","011010010010011000","010001100001010000","010001010010011000","011010011000000000");
		constant e_7 :pieces :=( "000000000000000000","000000000000000000","000011010010010011","000010001100001010","000011010010001010","000000000011010011");
		constant f_0 :pieces :=( "000000000000000000","000011010011000000","000010001010011000","000010100001010000","000010001010011000","000011010011000000");
		constant f_1 :pieces :=( "000000000000000000","000000011010011000","000011010001010000","000010001100010000","000011010001010000","000000011010011000");
		constant f_2 :pieces :=( "000011010011000000","000010001010011000","000010100001010000","000010001010011000","000011010011000000","000000000000000000");
		constant f_3 :pieces :=( "000000011010011000","000011010001010000","000010001100010000","000011010001010000","000000011010011000","000000000000000000");
		constant f_4 :pieces :=( "000000000000000000","011010010010011000","010001100001010000","011010001010011000","000011010011000000","000000000000000000");
		constant f_5 :pieces :=( "000000000000000000","000011010010010011","000010001100001010","000011010001010011","000000011010011000","000000000000000000");
		constant f_6 :pieces :=( "000000000000000000","000011010011000000","011010001010011000","010001100001010000","011010010010011000","000000000000000000");
		constant f_7 :pieces :=( "000000000000000000","000000011010011000","000011010001010011","000010001100001010","000011010010010011","000000000000000000");
		constant g_0 :pieces :=( "000000000000000000","000000000000000000","000011010010011000","000010100001010000","000010001001010000","000011010010011000");
		constant g_1 :pieces :=( "000000000000000000","000000000000000000","000011010010011000","000010001100010000","000010001001010000","000011010010011000");
		constant g_2 :pieces :=( "000011010010011000","000010001001010000","000010100001010000","000011010010011000","000000000000000000","000000000000000000");
		constant g_3 :pieces :=( "000011010010011000","000010001001010000","000010001100010000","000011010010011000","000000000000000000","000000000000000000");
		constant g_4 :pieces :=( "000000000000000000","011010010011000000","010001100010000000","010001001010000000","011010010011000000","000000000000000000");
		constant g_5 :pieces :=( "000000000000000000","000000011010010011","000000010100001010","000000010001001010","000000011010010011","000000000000000000");
		constant g_6 :pieces :=( "000000000000000000","011010010011000000","010001001010000000","010001100010000000","011010010011000000","000000000000000000");
		constant g_7 :pieces :=( "000000000000000000","000000011010010011","000000010001001010","000000010100001010","000000011010010011","000000000000000000");
		constant h_0 :pieces :=( "000000000000000000","000000000000000000","011010010011000000","010001100010011000","011010001001010000","000011010010011000");
		constant h_1 :pieces :=( "000000000000000000","000000000000000000","000000011010010011","000011010100001010","000010001001010011","000011010010011000");
		constant h_2 :pieces :=( "000011010010011000","011010001001010000","010001100010011000","011010010011000000","000000000000000000","000000000000000000");
		constant h_3 :pieces :=( "000011010010011000","000010001001010011","000011010100001010","000000011010010011","000000000000000000","000000000000000000");
		constant h_4 :pieces :=( "000011010011000000","011010001010000000","010001100010000000","010001010011000000","011010011000000000","000000000000000000");
		constant h_5 :pieces :=( "000000011010011000","000000010001010011","000000010100001010","000000011010001010","000000000011010011","000000000000000000");
		constant h_6 :pieces :=( "000000000000000000","011010011000000000","010001010011000000","010001100010000000","011010001010000000","000011010011000000");
		constant h_7 :pieces :=( "000000000000000000","000000000011010011","000000011010001010","000000010100001010","000000010001010011","000000011010011000");
		constant i_0 :pieces :=( "000011010011000000","000010001010000000","011010001010000000","010001100010000000","010001010011000000","011010011000000000");
		constant i_1 :pieces :=( "000000011010011000","000000010001010000","000000010001010011","000000010100001010","000000011010001010","000000000011010011");
		constant i_2 :pieces :=( "011010011000000000","010001010011000000","010001100010000000","011010001010000000","000010001010000000","000011010011000000");
		constant i_3 :pieces :=( "000000000011010011","000000011010001010","000000010100001010","000000010001010011","000000010001010000","000000011010011000");
		constant i_4 :pieces :=( "011010010011000000","010001001010010011","011010100001001010","000011010010010011","000000000000000000","000000000000000000");
		constant i_5 :pieces :=( "000000011010010011","011010010001001010","010001001100010011","011010010010011000","000000000000000000","000000000000000000");
		constant i_6 :pieces :=( "000000000000000000","000000000000000000","000011010010010011","011010100001001010","010001001010010011","011010010011000000");
		constant i_7 :pieces :=( "000000000000000000","000000000000000000","011010010010011000","010001001100010011","011010010001001010","000000011010010011");
		constant j_0 :pieces :=( "000000000000000000","000011010011000000","011010001010000000","010001100010000000","010001001010000000","011010010011000000");
		constant j_1 :pieces :=( "000000000000000000","000000011010011000","000000010001010011","000000010100001010","000000010001001010","000000011010010011");
		constant j_2 :pieces :=( "011010010011000000","010001001010000000","010001100010000000","011010001010000000","000011010011000000","000000000000000000");
		constant j_3 :pieces :=( "000000011010010011","000000010001001010","000000010100001010","000000010001010011","000000011010011000","000000000000000000");
		constant j_4 :pieces :=( "011010010011000000","010001001010011000","010001100001010000","011010010010011000","000000000000000000","000000000000000000");
		constant j_5 :pieces :=( "000000011010010011","000011010001001010","000010001100001010","000011010010010011","000000000000000000","000000000000000000");
		constant j_6 :pieces :=( "000000000000000000","000000000000000000","011010010010011000","010001100001010000","010001001010011000","011010010011000000");
		constant j_7 :pieces :=( "000000000000000000","000000000000000000","000011010010010011","000010001100001010","000011010001001010","000000011010010011");
		constant k_0 :pieces :=( "000000000000000000","011010010011000000","010001001010000000","011010100010000000","010001001010000000","011010010011000000");
		constant k_1 :pieces :=( "000000000000000000","000000011010010011","000000010001001010","000000010100010011","000000010001001010","000000011010010011");
		constant k_2 :pieces :=( "011010010011000000","010001001010000000","011010100010000000","010001001010000000","011010010011000000","000000000000000000");
		constant k_3 :pieces :=( "000000011010010011","000000010001001010","000000010100010011","000000010001001010","000000011010010011","000000000000000000");
		constant k_4 :pieces :=( "011010011010011000","010001010001010000","010001100001010000","011010010010011000","000000000000000000","000000000000000000");
		constant k_5 :pieces :=( "000011010011010011","000010001010001010","000010001100001010","000011010010010011","000000000000000000","000000000000000000");
		constant k_6 :pieces :=( "000000000000000000","000000000000000000","011010010010011000","010001100001010000","010001010001010000","011010011010011000");
		constant k_7 :pieces :=( "000000000000000000","000000000000000000","000011010010010011","000010001100001010","000010001010001010","000011010011010011");
		constant l_0 :pieces :=( "000000000000000000","000011010011000000","000010001010000000","011010100010011000","010001001001010000","011010010010011000");
		constant l_1 :pieces :=( "000000000000000000","000000011010011000","000000010001010000","000011010100010011","000010001001001010","000011010010010011");
		constant l_2 :pieces :=( "011010010010011000","010001001001010000","011010100010011000","000010001010000000","000011010011000000","000000000000000000");
		constant l_3 :pieces :=( "000011010010010011","000010001001001010","000011010100010011","000000010001010000","000000011010011000","000000000000000000");
		constant l_4 :pieces :=( "011010011000000000","010001010010011000","010001100001010000","010001010010011000","011010011000000000","000000000000000000");
		constant l_5 :pieces :=( "000000000011010011","000011010010001010","000010001100001010","000011010010001010","000000000011010011","000000000000000000");
		constant l_6 :pieces :=( "000000000000000000","011010011000000000","010001010010011000","010001100001010000","010001010010011000","011010011000000000");
		constant l_7 :pieces :=( "000000000000000000","000000000011010011","000011010010001010","000010001100001010","000011010010001010","000000000011010011");
		constant m_0 :pieces :=( "000011010011000000","000010001010000000","000010001010010011","000010100001001010","000011010010010011","000000000000000000");
		constant m_1 :pieces :=( "000000011010011000","000000010001010000","011010010001010000","010001001100010000","011010010010011000","000000000000000000");
		constant m_2 :pieces :=( "000000000000000000","000011010010010011","000010100001001010","000010001010010011","000010001010000000","000011010011000000");
		constant m_3 :pieces :=( "000000000000000000","011010010010011000","010001001100010000","011010010001010000","000000010001010000","000000011010011000");
		constant m_4 :pieces :=( "000000000000000000","000011010010010011","000010100001001010","000010001010010011","000010001010000000","000011010011000000");
		constant m_5 :pieces :=( "000000000000000000","011010010010011000","010001001100010000","011010010001010000","000000010001010000","000000011010011000");
		constant m_6 :pieces :=( "000011010011000000","000010001010000000","000010001010010011","000010100001001010","000011010010010011","000000000000000000");
		constant m_7 :pieces :=( "000000011010011000","000000010001010000","011010010001010000","010001001100010000","011010010010011000","000000000000000000");
		constant n_0 :pieces :=( "000000000000000000","011010010011000000","010001001010011000","011010100001010000","000011010001010000","000000011010011000");
		constant n_1 :pieces :=( "000000000000000000","000000011010010011","000011010001001010","000010001100010011","000010001010011000","000011010011000000");
		constant n_2 :pieces :=( "000000011010011000","000011010001010000","011010100001010000","010001001010011000","011010010011000000","000000000000000000");
		constant n_3 :pieces :=( "000011010011000000","000010001010011000","000010001100010011","000011010001001010","000000011010010011","000000000000000000");
		constant n_4 :pieces :=( "000000011010011000","000011010001010000","011010100001010000","010001001010011000","011010010011000000","000000000000000000");
		constant n_5 :pieces :=( "000011010011000000","000010001010011000","000010001100010011","000011010001001010","000000011010010011","000000000000000000");
		constant n_6 :pieces :=( "000000000000000000","011010010011000000","010001001010011000","011010100001010000","000011010001010000","000000011010011000");
		constant n_7 :pieces :=( "000000000000000000","000000011010010011","000011010001001010","000010001100010011","000010001010011000","000011010011000000");
		constant o_0 :pieces :=( "000000000000000000","011010011000000000","010001010010011000","010001100001010000","011010010001010000","000000011010011000");
		constant o_1 :pieces :=( "000000000000000000","000000000011010011","000011010010001010","000010001100001010","000010001010010011","000011010011000000");
		constant o_2 :pieces :=( "000000011010011000","011010010001010000","010001100001010000","010001010010011000","011010011000000000","000000000000000000");
		constant o_3 :pieces :=( "000011010011000000","000010001010010011","000010001100001010","000011010010001010","000000000011010011","000000000000000000");
		constant o_4 :pieces :=( "000011010010011000","000010001001010000","011010100010011000","010001001010000000","011010010011000000","000000000000000000");
		constant o_5 :pieces :=( "000011010010011000","000010001001010000","000011010100010011","000000010001001010","000000011010010011","000000000000000000");
		constant o_6 :pieces :=( "000000000000000000","011010010011000000","010001001010000000","011010100010011000","000010001001010000","000011010010011000");
		constant o_7 :pieces :=( "000000000000000000","000000011010010011","000000010001001010","000011010100010011","000010001001010000","000011010010011000");
		constant p_0 :pieces :=( "000000000000000000","011010011000000000","010001010010011000","010001100001010000","011010001010011000","000011010011000000");
		constant p_1 :pieces :=( "000000000000000000","000000000011010011","000011010010001010","000010001100001010","000011010001010011","000000011010011000");
		constant p_2 :pieces :=( "000011010011000000","011010001010011000","010001100001010000","010001010010011000","011010011000000000","000000000000000000");
		constant p_3 :pieces :=( "000000011010011000","000011010001010011","000010001100001010","000011010010001010","000000000011010011","000000000000000000");
		constant p_4 :pieces :=( "000011010010011000","011010001001010000","010001100010011000","011010001010000000","000011010011000000","000000000000000000");
		constant p_5 :pieces :=( "000011010010011000","000010001001010011","000011010100001010","000000010001010011","000000011010011000","000000000000000000");
		constant p_6 :pieces :=( "000000000000000000","000011010011000000","011010001010000000","010001100010011000","011010001001010000","000011010010011000");
		constant p_7 :pieces :=( "000000000000000000","000000011010011000","000000010001010011","000011010100001010","000010001001010011","000011010010011000");
		constant q_0 :pieces :=( "000000000000000000","000011010011000000","011010001010011000","010001100001010000","011010001010011000","000011010011000000");
		--constant q_1 :pieces :=( "000000000000000000","000000011010011000","000011010001010011","000010001100001010","000011010001010011","000000011010011000");
		--constant q_2 :pieces :=( "000011010011000000","011010001010011000","010001100001010000","011010001010011000","000011010011000000","000000000000000000");
		--constant q_3 :pieces :=( "000000011010011000","000011010001010011","000010001100001010","000011010001010011","000000011010011000","000000000000000000");
		--constant q_4 :pieces :=( "000011010011000000","011010001010011000","010001100001010000","011010001010011000","000011010011000000","000000000000000000");
		--constant q_5 :pieces :=( "000000011010011000","000011010001010011","000010001100001010","000011010001010011","000000011010011000","000000000000000000");
		--constant q_6 :pieces :=( "000000000000000000","000011010011000000","011010001010011000","010001100001010000","011010001010011000","000011010011000000");
		--constant q_7 :pieces :=(	"000000000000000000","000000011010011000","000011010001010011","000010001100001010","000011010001010011","000000011010011000");


begin	
--p <= (5 => ( 0|3|6|9|12|15|18|21|24|27|30|33=> '1' , others => '0') ,others =>( others=> '0') );   -- for test bench
--a <= "hello1";

-------------------------- registers -----------------------------
process (clk)
begin
	if (clk'event and clk='1') then
		state_reg <= state_next;
		sw2 <= sw2_next;
		sw1 <= sw1_next;
		load_reg <= load_next;
		rotate <= rotate_next;
		P <= P_next;
		formnex <= formnex_next;
		form <= form_next;
		dout_reg <= dout_next;
		M_reg <= M;
		opp <= opp_next;
		x_reg <= x_next;
		y_reg <= y_next;
		data_code_ch_reg <= data_code_ch_next;

	end if;

end process;

x_in <= to_integer( unsigned( din(117 downto 113) ) ) ;
y_in <= to_integer( unsigned( din(112 downto 108) ) ) ;
--------------------------- data out --------------------------
ok <= dout_reg;
load <= load_reg;
data_code_ch <= data_code_ch_reg;
-------------------------- states ------------------------------

process(data_code_ch_reg,state_reg,load_reg,sw1,sw2,rotate,form,formnex,dout_reg,data_rec,M_reg,P,opp,x_reg,y_reg,round,din,x_in,y_in,load_code)

variable r,z: integer := 0; 
variable a: integer := 0;
variable allow : std_logic := '1';
begin 
	P_next <= P; 
	load_next <= load_reg;
	sw1_next <= sw1;	
	sw2_next <= sw2;	
	state_next <= state_reg;
	rotate_next <= rotate;
	form_next <= form;
	formnex_next <= formnex; 
	dout_next <= dout_reg;
	M <= M_reg;
	x_next <= x_reg;
	y_next <= y_reg;
	opp_next <= opp;
	data_code_ch_next <= data_code_ch_reg;
	
	case state_reg is 
			when "00" => 
					data_code_ch_next <= '0';
					sw1_next <= '0';
					sw2_next <= '0';
					if(load_code = '1') then
						load_next <= '0';
					else
						load_next <= '1';
					end if;
					if(data_rec = '1') then
						data_code_ch_next <= '1';
						if (round = "01") then
							M <= q_0;
							sw1_next <= '0';
							sw2_next <= '1';
							x_next <= 4;
							y_next <= 3;
						state_next <= "10";
					elsif (round = "10") then --------- 1st round q selected
							M <= q_0;
							sw1_next <= '0';
							sw2_next <= '1';
							x_next <= 4;
							y_next <= 3;
						state_next <= "10";
												------------------------------- opponent_mapping -------------------------------
						for i in 0 to 5 loop 
							for j in 0 to 5 loop 
								if ( x_in - i > 2 and x_in -i < 15 and y_in - j > 2 and y_in - j < 15) then
									opp_next( x_in - i - 3 ) ( ( (y_in - j - 3) * 3)+2   downto ( ( (y_in -j-3) * 3) ) ) <= din( (107-18*i-3*j) downto (108-18*i-3*(j+1) ) );
								end if;		
							end loop;
						end loop;
			------------------------------ form and rotate selection -------------------------
					else 	
						state_next <= "01";
					------------------------------- opponent_mapping -------------------------------
						for i in 0 to 5 loop 
							for j in 0 to 5 loop 
								if ( x_in - i > 2 and x_in -i < 15 and y_in - j > 2 and y_in - j < 15) then
									opp_next( x_in - i - 3 ) ( ( (y_in - j - 3) * 3)+2   downto ( ( (y_in -j-3) * 3) ) ) <= din( (107-18*i-3*j) downto (108-18*i-3*(j+1) ) );
								end if;		
							end loop;
						end loop;
			------------------------------ form and rotate selection -------------------------
												-------- priority 2 : n
						if( form (13) = '0' and formnex (13) = '0') then
							if (rotate(0) = '0') then
								rotate_next(0) <= '1';
								M <= n_0;
							elsif (rotate(1) = '0') then
								rotate_next(1) <= '1';
								M <= n_1;
							elsif (rotate(2) = '0') then
								rotate_next(2) <= '1';	
								M <= n_2;
							elsif (rotate(3) = '0') then
								rotate_next(3) <= '1';
								M <= n_3;
							elsif (rotate(4) = '0') then
								rotate_next(4) <= '1';
								M <= n_4;
							elsif (rotate(5) = '0') then
								rotate_next(5) <= '1';
								M <= n_5;
							elsif (rotate(6) = '0') then
								M <= n_6;
								rotate_next(6) <= '1';
							elsif (rotate(7) = '0') then
								M <= n_7;
								rotate_next <= (others => '0');
								formnex_next(13) <= '1';
							end if;
											-------- priority 3 : p
						elsif( form (15) = '0' and formnex (15) = '0' ) then
							if (rotate(0) = '0') then
								M <= p_0;
								rotate_next(0) <= '1';
							elsif (rotate(1) = '0') then
								M <= p_1;
								rotate_next(1) <= '1';
							elsif (rotate(2) = '0') then
								M <= p_2;
								rotate_next(2) <= '1';
							elsif (rotate(3) = '0') then
								rotate_next(3) <= '1';
								M <= p_3;
							elsif (rotate(4) = '0') then
								M <= p_4;
								rotate_next(4) <= '1';
							elsif (rotate(5) = '0') then
								M <= p_5;
								rotate_next(5) <= '1';
							elsif (rotate(6) = '0') then
								M <= p_6;
								rotate_next(6) <= '1';
							elsif (rotate(7) = '0') then
								M <= p_7;
								rotate_next <= (others => '0');
								formnex_next(15) <= '1';
							end if;
										-------- priority 4 : i
						elsif( form (8) = '0' and formnex (8) = '0' ) then
							if (rotate(0) = '0') then
								M <= i_0;
								rotate_next(0) <= '1';
							elsif (rotate(1) = '0') then
								M <= i_1;
								rotate_next(1) <= '1';
							elsif (rotate(2) = '0') then
								M <= i_2;
								rotate_next(2) <= '1';
							elsif (rotate(3) = '0') then
								M <= i_3;
								rotate_next(3) <= '1';
							elsif (rotate(4) = '0') then
								M <= i_4;
								rotate_next(4) <= '1';
							elsif (rotate(5) = '0') then
								M <= i_5;
								rotate_next(5) <= '1';
							elsif (rotate(6) = '0') then
								M <= i_6;
								rotate_next(6) <= '1';
							elsif (rotate(7) = '0') then
								M <= i_7;
								rotate_next <= (others => '0');
								formnex_next(8) <= '1';
							end if;
										-------- priority 5 : o
						elsif( form (14) = '0' and formnex (14) = '0') then
							if (rotate(0) = '0') then
								M <= o_0;
								rotate_next(0) <= '1';
							elsif (rotate(1) = '0') then
								M <= o_1;
								rotate_next(1) <= '1';
							elsif (rotate(2) = '0') then
								M <= o_2;
								rotate_next(2) <= '1';
							elsif (rotate(3) = '0') then
								M <= o_3;
								rotate_next(3) <= '1';
							elsif (rotate(4) = '0') then
								M <= o_4;
								rotate_next(4) <= '1';
							elsif (rotate(5) = '0') then
								M <= o_5;
								rotate_next(5) <= '1';
							elsif (rotate(6) = '0') then
								M <= o_6;
								rotate_next(6) <= '1';
							elsif (rotate(7) = '0') then
								M <= o_7;
								rotate_next <= (others => '0');
								formnex_next(14) <= '1';
							end if;
									-------- priority 6 : l
						elsif( form (11) = '0' and formnex (11) = '0') then
							if (rotate(0) = '0') then
								M <= l_0;
								rotate_next(0) <= '1';
							elsif (rotate(1) = '0') then
								M <= l_1;
								rotate_next(1) <= '1';
							elsif (rotate(2) = '0') then
								M <= l_2;
								rotate_next(2) <= '1';
							elsif (rotate(3) = '0') then
								M <= l_3;
								rotate_next(3) <= '1';
							elsif (rotate(4) = '0') then
								M <= l_4;
								rotate_next(4) <= '1';
							elsif (rotate(5) = '0') then
								M <= l_5;
								rotate_next(5) <= '1';
							elsif (rotate(6) = '0') then
								M <= l_6;
								rotate_next(6) <= '1';
							elsif (rotate(7) = '0') then
								M <= l_7;
								rotate_next <= (others => '0');
								formnex_next(11) <= '1';
							end if;
									-------- priority 7 : j
						elsif( form (9) = '0' and formnex (9) = '0') then
							if (rotate(0) = '0') then
								M <= j_0;
								rotate_next(0) <= '1';
							elsif (rotate(1) = '0') then
								M <= j_1;
								rotate_next(1) <= '1';
							elsif (rotate(2) = '0') then
								M <= j_2;
								rotate_next(2) <= '1';
							elsif (rotate(3) = '0') then
								M <= j_3;
								rotate_next(3) <= '1';
							elsif (rotate(4) = '0') then
								M <= j_4;
								rotate_next(4) <= '1';
							elsif (rotate(5) = '0') then
								M <= j_5;
								rotate_next(5) <= '1';
							elsif (rotate(6) = '0') then
								M <= j_6;
								rotate_next(6) <= '1';
							elsif (rotate(7) = '0') then
								M <= j_7;
								formnex_next(9) <= '1';
								rotate_next <= (others => '0');
							end if;
									-------- priority 8 : k
						elsif( form (10) = '0' and formnex (10) = '0') then
							if (rotate(0) = '0') then
								M <= k_0;
								rotate_next(0) <= '1';
							elsif (rotate(1) = '0') then
								M <= k_1;
								rotate_next(1) <= '1';
							elsif (rotate(2) = '0') then
								M <= k_2;
								rotate_next(2) <= '1';
							elsif (rotate(3) = '0') then
								M <= k_3;
								rotate_next(3) <= '1';
							elsif (rotate(4) = '0') then
								M <= k_4;
								rotate_next(4) <= '1';
							elsif (rotate(5) = '0') then
								M <= k_5;
								rotate_next(5) <= '1';
							elsif (rotate(6) = '0') then
								M <= k_6;
								rotate_next(6) <= '1';
							elsif (rotate(7) = '0') then
								M <= k_7;
								formnex_next(10) <= '1';
								rotate_next <= (others => '0');
							end if;
									-------- priority 9 : m
						elsif( form (12) = '0' and formnex (12) = '0') then
							if (rotate(0) = '0') then
								M <= m_0;
								rotate_next(0) <= '1';
							elsif (rotate(1) = '0') then
								M <= m_1;
								rotate_next(1) <= '1';
							elsif (rotate(2) = '0') then
								M <= m_2;
								rotate_next(2) <= '1';
							elsif (rotate(3) = '0') then
								M <= m_3;
								rotate_next(3) <= '1';
							elsif (rotate(4) = '0') then
								M <= m_4;
								rotate_next(4) <= '1';
							elsif (rotate(5) = '0') then
								M <= m_5;
								rotate_next(5) <= '1';
							elsif (rotate(6) = '0') then
								M <= m_6;
								rotate_next(6) <= '1';
							elsif (rotate(7) = '0') then
								M <= m_7;
								formnex_next(12) <= '1';
								rotate_next <= (others => '0');
							end if;
									-------- priority 10 : h
						elsif( form (7) = '0' and formnex (7) = '0') then
							if (rotate(0) = '0') then
								M <= h_0;
								rotate_next(0) <= '1';
							elsif (rotate(1) = '0') then
								M <= h_1;
								rotate_next(1) <= '1';
							elsif (rotate(2) = '0') then
								M <= h_2;
								rotate_next(2) <= '1';
							elsif (rotate(3) = '0') then
								M <= h_3;
								rotate_next(3) <= '1';
							elsif (rotate(4) = '0') then
								M <= h_4;
								rotate_next(4) <= '1';
							elsif (rotate(5) = '0') then
								M <= h_5;
								rotate_next(5) <= '1';
							elsif (rotate(6) = '0') then
								M <= h_6;
								rotate_next(6) <= '1';
							elsif (rotate(7) = '0') then
								M <= h_7;
								formnex_next(7) <= '1';
								rotate_next <= (others => '0');
							end if;
									-------- priority 11 : f
						elsif( form (5) = '0' and formnex (5) = '0') then
							if (rotate(0) = '0') then
								M <= f_0;
								rotate_next(0) <= '1';
							elsif (rotate(1) = '0') then
								M <= f_1;
								rotate_next(1) <= '1';
							elsif (rotate(2) = '0') then
								M <= f_2;
								rotate_next(2) <= '1';
							elsif (rotate(3) = '0') then
								M <= f_3;
								rotate_next(3) <= '1';
							elsif (rotate(4) = '0') then
								M <= f_4;
								rotate_next(4) <= '1';
							elsif (rotate(5) = '0') then
								M <= f_5;
								rotate_next(5) <= '1';
							elsif (rotate(6) = '0') then
								M <= f_6;
								rotate_next(6) <= '1';
							elsif (rotate(7) = '0') then
								M <= f_7;
								formnex_next(5) <= '1';
								rotate_next <= (others => '0');
							end if;
									-------- priority 12 : e
						elsif( form (4) = '0' and formnex (4) = '0') then
							if (rotate(0) = '0') then
								M <= e_0;
								rotate_next(0) <= '1';
							elsif (rotate(1) = '0') then
								M <= e_1;
								rotate_next(1) <= '1';
							elsif (rotate(2) = '0') then
								M <= e_2;
								rotate_next(2) <= '1';
							elsif (rotate(3) = '0') then
								M <= e_3;
								rotate_next(3) <= '1';
							elsif (rotate(4) = '0') then
								M <= e_4;
								rotate_next(4) <= '1';
							elsif (rotate(5) = '0') then
								M <= e_5;
								rotate_next(5) <= '1';
							elsif (rotate(6) = '0') then
								M <= e_6;
								rotate_next(6) <= '1';
							elsif (rotate(7) = '0') then
								M <= e_7;
								formnex_next(4) <= '1';
								rotate_next <= (others => '0');
							end if;
									-------- priority 13 : g
						elsif( form (6) = '0' and formnex (6) = '0') then
							if (rotate(0) = '0') then
								M <= g_0;
								rotate_next(0) <= '1';
							elsif (rotate(1) = '0') then
								M <= g_1;
								rotate_next(1) <= '1';
							elsif (rotate(2) = '0') then
								M <= g_2;
								rotate_next(2) <= '1';
							elsif (rotate(3) = '0') then
								M <= g_3;
								rotate_next(3) <= '1';
							elsif (rotate(4) = '0') then
								M <= g_4;
								rotate_next(4) <= '1';
							elsif (rotate(5) = '0') then
								M <= g_5;
								rotate_next(5) <= '1';
							elsif (rotate(6) = '0') then
								M <= g_6;
								rotate_next(6) <= '1';
							elsif (rotate(7) = '0') then
								M <= g_7;
								formnex_next(6) <= '1';
								rotate_next <= (others => '0');
							end if;
									-------- priority 14 : d
						elsif( form (3) = '0' and formnex (3) = '0') then
							if (rotate(0) = '0') then
								M <= d_0;
								rotate_next(0) <= '1';
							elsif (rotate(1) = '0') then
								M <= d_1;
								rotate_next(1) <= '1';
							elsif (rotate(2) = '0') then
								M <= d_2;
								rotate_next(2) <= '1';
							elsif (rotate(3) = '0') then
								M <= d_3;
								rotate_next(3) <= '1';
							elsif (rotate(4) = '0') then
								M <= d_4;
								rotate_next(4) <= '1';
							elsif (rotate(5) = '0') then
								M <= d_5;
								rotate_next(5) <= '1';
							elsif (rotate(6) = '0') then
								M <= d_6;
								rotate_next(6) <= '1';
							elsif (rotate(7) = '0') then
								M <= d_7;
								formnex_next(3) <= '1';
								rotate_next <= (others => '0');
							end if;
									-------- priority 15 : c
						elsif( form (2) = '0' and formnex (2) = '0') then
							if (rotate(0) = '0') then
								M <= c_0;
								rotate_next(0) <= '1';
							elsif (rotate(1) = '0') then
								M <= c_1;
								rotate_next(1) <= '1';
							elsif (rotate(2) = '0') then
								M <= c_2;
								rotate_next(2) <= '1';
							elsif (rotate(3) = '0') then
								M <= c_3;
								rotate_next(3) <= '1';
							elsif (rotate(4) = '0') then
								M <= c_4;
								rotate_next(4) <= '1';
							elsif (rotate(5) = '0') then
								M <= c_5;
								rotate_next(5) <= '1';
							elsif (rotate(6) = '0') then
								M <= c_6;
								rotate_next(6) <= '1';
							elsif (rotate(7) = '0') then
								M <= c_7;
								formnex_next(2) <= '1';
								rotate_next <= (others => '0');
							end if;
									-------- priority 16 : b
						elsif( form (1) = '0' and formnex (1) = '0') then
							if (rotate(0) = '0') then
								M <= b_0;
								rotate_next(0) <= '1';
							elsif (rotate(1) = '0') then
								M <= b_1;
								rotate_next(1) <= '1';
							elsif (rotate(2) = '0') then
								M <= b_2;
								rotate_next(2) <= '1';
							elsif (rotate(3) = '0') then
								M <= b_3;
								rotate_next(3) <= '1';
							elsif (rotate(4) = '0') then
								M <= b_4;
								rotate_next(4) <= '1';
							elsif (rotate(5) = '0') then
								M <= b_5;
								rotate_next(5) <= '1';
							elsif (rotate(6) = '0') then
								M <= b_6;
								rotate_next(6) <= '1';
							elsif (rotate(7) = '0') then
								M <= b_7;
								formnex_next(1) <= '1';
								rotate_next <= (others => '0');
							end if;
									-------- priority 17 : a
						elsif( form (0) = '0' and formnex (13) = '0') then
							if (rotate(0) = '0') then
								M <= a_0;
								rotate_next(0) <= '1';
							elsif (rotate(1) = '0') then
								M <= a_1;
								rotate_next(1) <= '1';
							elsif (rotate(2) = '0') then
								M <= a_2;
								rotate_next(2) <= '1';
							elsif (rotate(3) = '0') then
								M <= a_3;
								rotate_next(3) <= '1';
							elsif (rotate(4) = '0') then
								M <= a_4;
								rotate_next(4) <= '1';
							elsif (rotate(5) = '0') then
								M <= a_5;
								rotate_next(5) <= '1';
							elsif (rotate(6) = '0') then
								M <= a_6;
								rotate_next(6) <= '1';
							elsif (rotate(7) = '0') then
								M <= a_7;
								formnex_next(0) <= '1';
								rotate_next <= (others => '0');
							end if;
						end if;
					  end if;
					else 
						state_next <= "00";
					end if;
		when "01" =>  			
								-------------------------- check the conditions for puting a piece ---------------------------
						state_next <= "10";
	--for x in 0 to 17 loop
		--for y in 0 to 17 loop
		--	if ( y >= 15 or x >=15) then
		--		exit;
		--	end if;
			for i in 0 to 5 loop
				for j in 0 to 5 loop
					allow := '1';
					r := i+x_reg;
					z := j+y_reg;
					if (x_reg < 3) then
						if( (i < (3 - x_reg)) and ( (M_reg(i)( ((j*3)+2) downto (j*3) ) = "001") or  (M_reg(i)( ((j*3)+2) downto (j*3) ) = "100")) ) then
							sw1_next <= '1';
							exit;
						end if;
						if ( i < (3 - x_reg) ) then
							allow := '0';
						end if;
						r := i+ x_reg -3;
					end if;
				if (y_reg < 3) then
						if( (j < (3-y_reg)) and ( (M_reg(i)( ((j*3)+2) downto (j*3) ) = "001") or  (M_reg(i)( ((j*3)+2) downto (j*3) ) = "100")) ) then
							sw1_next <= '1';
							exit;
						end if;
						if ( j < (3-y_reg) ) then
							allow := '0';
						end if;
 						z := j+y_reg-3;	 
					end if;
					if (x_reg > 9 and x_reg < 15) then
						if( (i > (14-x_reg)) and ( (M_reg(i)( ((j*3)+2) downto (j*3) ) = "001") or  (M_reg(i)( ((j*3)+2) downto (j*3) ) = "100")) ) then
							sw1_next <= '1';
							exit;
						end if;	 
						if ( i > (14-x_reg) ) then
							allow := '0';
						end if;
					end if;
					if (y_reg > 9 and y_reg < 15) then
						if( (j > (14-y_reg)) and ( (M_reg(i)( ((j*3)+2) downto (j*3) ) = "001") or  (M_reg(i)( ((j*3)+2) downto (j*3) ) = "100")) ) then
							sw1_next <= '1';
							exit;
						end if;	 
						if ( j > (14-y_reg) )then
							allow := '0';
						end if;
					end if;
					if (allow = '1') then
						if( (P(r)( ((z*3)+2) downto (z*3) ) = "001") and  ( (M_reg(i)( ((j*3)+2) downto (j*3) ) = "100") or (M_reg(i)( ((j*3)+2) downto (j*3) ) = "001")) ) then
								sw1_next <= '1';
								exit;
							end if;	 		
						if (M_reg(i)(j*3) = '0' and M_reg(i)((j*3)+1) = '1' and M_reg(i)((j*3)+2) = '0' and P(r)(z*3) = '1' and P(r)((z*3)+1) = '0' and P(r)((z*3)+2) = '0' ) then 
							sw1_next <= '1';
							exit ;
						end if;
						if( (opp(r)( ((z*3)+2) downto (z*3) ) = "001") and  ( (M_reg(i)( ((j*3)+2) downto (j*3) ) = "100") or (M_reg(i)( ((j*3)+2) downto (j*3) ) = "001")) ) then
								sw1_next <= '1';
								exit;
							end if;	
						if (M_reg(i)(j*3) = '1' and M_reg(i)((j*3)+1) = '1' and M_reg(i)((j*3)+2) = '0' and P(r)(z*3) = '1' and P(r)((z*3)+1) = '0' and P(r)((z*3)+2) = '0' ) then 
							sw2_next <= '1';
						end if;
					end if;	
				end loop;
			end loop;
	--	end loop;
	--end loop;
	when "10" =>
				if(sw2 = '1' and sw1 = '0') then
					dout_next <=(std_logic_vector(to_unsigned((x_reg+5),5)) & std_logic_vector(to_unsigned((y_reg+5),5)) & M_reg(5)(17 downto 0) 
					& M_reg(4)(17 downto 0) & M_reg(3)(17 downto 0) & M_reg(2)(17 downto 0) & M_reg(1)(17 downto 0) & M_reg(0)(17 downto 0));
					if (M_reg = n_0 or M_reg = n_1 or M_reg = n_2 or M_reg = n_3 or M_reg = n_4 or M_reg = n_5 or M_reg = n_6 or M_reg = n_7)	then 
						form_next(13) <= '1';
					elsif (M_reg = p_0 or M_reg = p_1 or M_reg = p_2 or M_reg = p_3 or M_reg = p_4 or M_reg = p_5 or M_reg = p_6 or M_reg = p_7)	then 
						form_next(15) <= '1';
					elsif (M_reg = i_0 or M_reg = i_1 or M_reg = i_2 or M_reg = i_3 or M_reg = i_4 or M_reg = i_5 or M_reg = i_6 or M_reg = i_7)	then 
						form_next(8) <= '1';
					elsif (M_reg = o_0 or M_reg = o_1 or M_reg = o_2 or M_reg = o_3 or M_reg = o_4 or M_reg = o_5 or M_reg = o_6 or M_reg = o_7)	then 
						form_next(14) <= '1';
					elsif (M_reg = l_0 or M_reg = l_1 or M_reg = l_2 or M_reg = l_3 or M_reg = l_4 or M_reg = l_5 or M_reg = l_6 or M_reg = l_7)	then 
						form_next(11) <= '1';
					elsif (M_reg = j_0 or M_reg = j_1 or M_reg = j_2 or M_reg = j_3 or M_reg = j_4 or M_reg = j_5 or M_reg = j_6 or M_reg = j_7)	then 
						form_next(9) <= '1';
					elsif (M_reg = k_0 or M_reg = k_1 or M_reg = k_2 or M_reg = k_3 or M_reg = k_4 or M_reg = k_5 or M_reg = k_6 or M_reg = k_7)	then 
						form_next(10) <= '1';
					elsif (M_reg = m_0 or M_reg = m_1 or M_reg = m_2 or M_reg = m_3 or M_reg = m_4 or M_reg = m_5 or M_reg = m_6 or M_reg = m_7)	then 
						form_next(12) <= '1';
					elsif (M_reg = h_0 or M_reg = h_1 or M_reg = h_2 or M_reg = h_3 or M_reg = h_4 or M_reg = h_5 or M_reg = h_6 or M_reg = h_7)	then 
						form_next(7) <= '1';
					elsif (M_reg = f_0 or M_reg = f_1 or M_reg = f_2 or M_reg = f_3 or M_reg = f_4 or M_reg = f_5 or M_reg = f_6 or M_reg = f_7)	then 
						form_next(5) <= '1';
					elsif (M_reg = e_0 or M_reg = e_1 or M_reg = e_2 or M_reg = e_3 or M_reg = e_4 or M_reg = e_5 or M_reg = e_6 or M_reg = e_7)	then 
						form_next(4) <= '1';
					elsif (M_reg = g_0 or M_reg = g_1 or M_reg = g_2 or M_reg = g_3 or M_reg = g_4 or M_reg = g_5 or M_reg = g_6 or M_reg = g_7)	then 
						form_next(6) <= '1';
					elsif (M_reg = d_0 or M_reg = d_1 or M_reg = d_2 or M_reg = d_3 or M_reg = d_4 or M_reg = d_5 or M_reg = d_6 or M_reg = d_7)	then 
						form_next(3) <= '1';
					elsif (M_reg = c_0 or M_reg = c_1 or M_reg = c_2 or M_reg = c_3 or M_reg = c_4 or M_reg = c_5 or M_reg = c_6 or M_reg = c_7)	then 
						form_next(2) <= '1';
					elsif (M_reg = b_0 or M_reg = b_1 or M_reg = b_2 or M_reg = b_3 or M_reg = b_4 or M_reg = b_5 or M_reg = b_6 or M_reg = b_7)	then 
						form_next(1) <= '1';
					elsif (M_reg = a_0 or M_reg = a_1 or M_reg = a_2 or M_reg = a_3 or M_reg = a_4 or M_reg = a_5 or M_reg = a_6 or M_reg = a_7)	then 
						form_next(0) <= '1';
					end if;				
					state_next <= "11";
					rotate_next <= (others => '0');
				end if;	
				if(	y_reg < 13 ) then 
					y_next <= y_reg+1;
					state_next <= "01";
				elsif ( x_reg < 13 ) then 
					x_next <= x_reg+1;
					y_next <= 0;
					state_next <= "01";
				else 
					x_next <= 0;
					y_next <= 0;
					state_next <= "00";	
				end if;
	when "11" =>
					load_next <= '1';
										--------------- our map ------------------
					for i in 0 to 5 loop 
						for j in 0 to 17 loop 
							if ( (x_reg+i) > 2 and (x_reg+i) < 15 and (y_reg * 3 + j) > 8 and (y_reg * 3 + j) < 45) then 
								P_next( x_reg + i - 3 ) ( y_reg * 3 + j - 9 ) <= dout_reg( 18*i+j );
							end if;		
						end loop;
					end loop;	
							-----------------------------------------------
				formnex_next <= form;
				state_next <= "00";
				x_next <= 0;
				y_next <= 0;
--	when "100" =>
--					--------------- delay for loading data------------
--				start_next <= '1';
--				load_next <= '0';
--				state_next <= "101";
--		when "101" =>
--						---------- delay for sending data ------------
--				state_next <= "000";
--	when others =>
--				state_next <= "000";
	end case;	
end process;

end failure;



--architecture test_bench of code is
--
--  -- Component Declaration
--Component x  port (
--ok : out std_logic_vector(117 downto 0);
--opponent : in std_logic_vector(431 downto 0);
--clk : in std_logic);
--end component;
-- 
--for g:x use Entity work.code(failure);
--
--signal ok1 : std_logic_vector(117 downto 0) ;
--signal clk1 : std_logic := '0';
--signal opponent1 : std_logic_vector(431 downto 0):= (1 => '1' , others => '0');
--begin
--
---- Component Instantiation
--  g: x PORT MAP(ok1,opponent1,clk1);
--
--    opponent1 <= (1 => '1' , others => '0') after 1 ns;
--		clk1 <= '1' after 3 ns,'0' after 4 ns,'1' after 5 ns,'0' after 6 ns,'1' after 7 ns,
--						'0' after 8 ns,'1' after 9 ns,'0' after 10 ns,'1' after 11 ns,'0' after 12 ns,'1' after 13 ns;
--
--end test_bench;
--
--
--

