library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std.All;

-------------------------------
---- Uncomment the following library declaration if instantiating
entity program is
    Port ( datain : in std_logic_vector(31 downto 0);
				  data_decoded : out std_logic_vector (117 downto 0);
					min_max_out : out unsigned (15 downto 0)
);
end program;
-------------------------------------
architecture Gate_level of program is

		type MATRIX is array(5 downto 0) of std_logic_vector(17 downto 0);
		type MIX is array(16 downto 0) of unsigned(15 downto 0);

		signal sampler : MATRIX := (others=>(others=>'0'));
		signal X_ini,Y_ini : unsigned(7 downto 0);
		signal X_ini_before,Y_ini_before : unsigned(7 downto 0);
		signal format : unsigned (7 downto 0);
		signal rotate : unsigned (7 downto 0);
		signal alaki : unsigned (5 downto 0);

		constant mix_array : MIX := (others=>(others=>'0'));

begin

		rotate <= 							"00000111"	when (datain(7 downto 0) = "00110111") else
									"00000110"	when (datain(7 downto 0) = "00110110") else
									"00000101"	when (datain(7 downto 0) = "00110101") else
									"00000100"	when (datain(7 downto 0) = "00110100") else
									"00000011"	when (datain(7 downto 0) = "00110011") else
									"00000010"	when (datain(7 downto 0) = "00110010") else
									"00000001"	when (datain(7 downto 0) = "00110001") else
									"00000000" ;


		format <= unsigned(datain(15 downto 8));

		X_ini_before <=	"00000011" when (datain(31 downto 24) = "01100011") else 
									"00000100" when (datain(31 downto 24) = "01100010") else
									"00000101" when (datain(31 downto 24) = "01100001") else
									"00000110"	when (datain(31 downto 24) = "00111001") else
									"00000111"	when (datain(31 downto 24) = "00111000") else
									"00001000"	when (datain(31 downto 24) = "00110111") else
									"00001001"	when (datain(31 downto 24) = "00110110") else
									"00001010"	when (datain(31 downto 24) = "00110101") else
									"00001011"	when (datain(31 downto 24) = "00110100") else
									"00001100"	when (datain(31 downto 24) = "00110011") else
									"00001101"	when (datain(31 downto 24) = "00110010") else
									"00001110"	when (datain(31 downto 24) = "00110001") else
									"00000000" ;

		X_ini <= X_ini_before +3	when (rotate = 0 or rotate = 2 or rotate = 4 or rotate = 6) else --rotate = 0|2|4|6
						X_ini_before +2;	--when (rotate = 1  or rotate = 3 or rotate = 5 or rotate = 7); --rotate = 1|3|5|7

		Y_ini_before <=	"00000011" when (datain(23 downto 16) = "01100011") else 
									"00000100" when (datain(23 downto 16) = "01100010") else
									"00000101" when (datain(23 downto 16) = "01100001") else
									"00000110"	when (datain(23 downto 16) = "00111001") else
									"00000111"	when (datain(23 downto 16) = "00111000") else
									"00001000"	when (datain(23 downto 16) = "00110111") else
									"00001001"	when (datain(23 downto 16) = "00110110") else
									"00001010"	when (datain(23 downto 16) = "00110101") else
									"00001011"	when (datain(23 downto 16) = "00110100") else
									"00001100"	when (datain(23 downto 16) = "00110011") else
									"00001101"	when (datain(23 downto 16) = "00110010") else
									"00001110"	when (datain(23 downto 16) = "00110001") else
									"00000000" ;
		Y_ini <= Y_ini_before +2	when (rotate = 0 or rotate = 1  or rotate = 6 or rotate = 7) else --rotate = 0|1|6|7
						Y_ini_before +3 ;--	when (rotate = 2 or rotate = 3 or rotate = 4 or rotate = 5);  --rotate = 2|3|4|5						


		sampler <=		( "000000000000000000","000000000000000000","000011010011000000","000010100010000000","000011010011000000","000000000000000000")	when  (format = 97 and rotate = 0) else
( "000000000000000000","000000000000000000","000000011010011000","000000010100010000","000000011010011000","000000000000000000")	when  (format = 97 and rotate = 1) else
( "000000000000000000","000011010011000000","000010100010000000","000011010011000000","000000000000000000","000000000000000000")	when  (format = 97 and rotate = 2) else
( "000000000000000000","000000011010011000","000000010100010000","000000011010011000","000000000000000000","000000000000000000")	when  (format = 97 and rotate = 3) else
( "000000000000000000","000011010011000000","000010100010000000","000011010011000000","000000000000000000","000000000000000000")	when  (format = 97 and rotate = 4) else
( "000000000000000000","000000011010011000","000000010100010000","000000011010011000","000000000000000000","000000000000000000")	when  (format = 97 and rotate = 5) else
( "000000000000000000","000000000000000000","000011010011000000","000010100010000000","000011010011000000","000000000000000000")	when  (format = 97 and rotate = 6) else
( "000000000000000000","000000000000000000","000000011010011000","000000010100010000","000000011010011000","000000000000000000")	when  (format = 97 and rotate = 7) else
( "000000000000000000","000000000000000000","000011010011000000","000010100010000000","000010001010000000","000011010011000000")	when  (format = 98 and rotate = 0) else
( "000000000000000000","000000000000000000","000000011010011000","000000010100010000","000000010001010000","000000011010011000")	when  (format = 98 and rotate = 1) else
( "000011010011000000","000010001010000000","000010100010000000","000011010011000000","000000000000000000","000000000000000000")	when  (format = 98 and rotate = 2) else
( "000000011010011000","000000010001010000","000000010100010000","000000011010011000","000000000000000000","000000000000000000")	when  (format = 98 and rotate = 3) else
( "000000000000000000","011010010011000000","010001100010000000","011010010011000000","000000000000000000","000000000000000000")	when  (format = 98 and rotate = 4) else
( "000000000000000000","000000011010010011","000000010100001010","000000011010010011","000000000000000000","000000000000000000")	when  (format = 98 and rotate = 5) else
( "000000000000000000","000000000000000000","011010010011000000","010001100010000000","011010010011000000","000000000000000000")	when  (format = 98 and rotate = 6) else
( "000000000000000000","000000000000000000","000000011010010011","000000010100001010","000000011010010011","000000000000000000")	when  (format = 98 and rotate = 7) else
( "000000000000000000","000011010011000000","000010001010000000","000010100010000000","000010001010000000","000011010011000000")	when  (format = 99 and rotate = 0) else
( "000000000000000000","000000011010011000","000000010001010000","000000010100010000","000000010001010000","000000011010011000")	when  (format = 99 and rotate = 1) else
( "000011010011000000","000010001010000000","000010100010000000","000010001010000000","000011010011000000","000000000000000000")	when  (format = 99 and rotate = 2) else
( "000000011010011000","000000010001010000","000000010100010000","000000010001010000","000000011010011000","000000000000000000")	when  (format = 99 and rotate = 3) else
( "000000000000000000","011010010010011000","010001100001010000","011010010010011000","000000000000000000","000000000000000000")	when  (format = 99 and rotate = 4) else
( "000000000000000000","000011010010010011","000010001100001010","000011010010010011","000000000000000000","000000000000000000")	when  (format = 99 and rotate = 5) else
( "000000000000000000","000000000000000000","011010010010011000","010001100001010000","011010010010011000","000000000000000000")	when  (format = 99 and rotate = 6) else
( "000000000000000000","000000000000000000","000011010010010011","000010001100001010","000011010010010011","000000000000000000")	when  (format = 99 and rotate = 7) else
( "000000000000000000","000011010011000000","000010001010011000","000010100001010000","000011010010011000","000000000000000000")	when  (format = 100 and rotate = 0) else
( "000000000000000000","000000011010011000","000011010001010000","000010001100010000","000011010010011000","000000000000000000")	when  (format = 100 and rotate = 1) else
( "000000000000000000","000011010010011000","000010100001010000","000010001010011000","000011010011000000","000000000000000000")	when  (format = 100 and rotate = 2) else
( "000000000000000000","000011010010011000","000010001100010000","000011010001010000","000000011010011000","000000000000000000")	when  (format = 100 and rotate = 3) else
( "000000000000000000","000011010010011000","000010100001010000","000010001010011000","000011010011000000","000000000000000000")	when  (format = 100 and rotate = 4) else
( "000000000000000000","000011010010011000","000010001100010000","000011010001010000","000000011010011000","000000000000000000")	when  (format = 100 and rotate = 5) else
( "000000000000000000","000011010011000000","000010001010011000","000010100001010000","000011010010011000","000000000000000000")	when  (format = 100 and rotate = 6) else
( "000000000000000000","000000011010011000","000011010001010000","000010001100010000","000011010010011000","000000000000000000")	when  (format = 100 and rotate = 7) else
( "000000000000000000","000011010011000000","000010001010000000","011010100010000000","010001001010000000","011010010011000000")	when  (format = 101 and rotate = 0) else
( "000000000000000000","000000011010011000","000000010001010000","000000010100010011","000000010001001010","000000011010010011")	when  (format = 101 and rotate = 1) else
( "011010010011000000","010001001010000000","011010100010000000","000010001010000000","000011010011000000","000000000000000000")	when  (format = 101 and rotate = 2) else
( "000000011010010011","000000010001001010","000000010100010011","000000010001010000","000000011010011000","000000000000000000")	when  (format = 101 and rotate = 3) else
( "011010011000000000","010001010010011000","010001100001010000","011010010010011000","000000000000000000","000000000000000000")	when  (format = 101 and rotate = 4) else
( "000000000011010011","000011010010001010","000010001100001010","000011010010010011","000000000000000000","000000000000000000")	when  (format = 101 and rotate = 5) else
( "000000000000000000","000000000000000000","011010010010011000","010001100001010000","010001010010011000","011010011000000000")	when  (format = 101 and rotate = 6) else
( "000000000000000000","000000000000000000","000011010010010011","000010001100001010","000011010010001010","000000000011010011")	when  (format = 101 and rotate = 7) else
( "000000000000000000","000011010011000000","000010001010011000","000010100001010000","000010001010011000","000011010011000000")	when  (format = 102 and rotate = 0) else
( "000000000000000000","000000011010011000","000011010001010000","000010001100010000","000011010001010000","000000011010011000")	when  (format = 102 and rotate = 1) else
( "000011010011000000","000010001010011000","000010100001010000","000010001010011000","000011010011000000","000000000000000000")	when  (format = 102 and rotate = 2) else
( "000000011010011000","000011010001010000","000010001100010000","000011010001010000","000000011010011000","000000000000000000")	when  (format = 102 and rotate = 3) else
( "000000000000000000","011010010010011000","010001100001010000","011010001010011000","000011010011000000","000000000000000000")	when  (format = 102 and rotate = 4) else
( "000000000000000000","000011010010010011","000010001100001010","000011010001010011","000000011010011000","000000000000000000")	when  (format = 102 and rotate = 5) else
( "000000000000000000","000011010011000000","011010001010011000","010001100001010000","011010010010011000","000000000000000000")	when  (format = 102 and rotate = 6) else
( "000000000000000000","000000011010011000","000011010001010011","000010001100001010","000011010010010011","000000000000000000")	when  (format = 102 and rotate = 7) else
( "000000000000000000","000000000000000000","000011010010011000","000010100001010000","000010001001010000","000011010010011000")	when  (format = 103 and rotate = 0) else
( "000000000000000000","000000000000000000","000011010010011000","000010001100010000","000010001001010000","000011010010011000")	when  (format = 103 and rotate = 1) else
( "000011010010011000","000010001001010000","000010100001010000","000011010010011000","000000000000000000","000000000000000000")	when  (format = 103 and rotate = 2) else
( "000011010010011000","000010001001010000","000010001100010000","000011010010011000","000000000000000000","000000000000000000")	when  (format = 103 and rotate = 3) else
( "000000000000000000","011010010011000000","010001100010000000","010001001010000000","011010010011000000","000000000000000000")	when  (format = 103 and rotate = 4) else
( "000000000000000000","000000011010010011","000000010100001010","000000010001001010","000000011010010011","000000000000000000")	when  (format = 103 and rotate = 5) else
( "000000000000000000","011010010011000000","010001001010000000","010001100010000000","011010010011000000","000000000000000000")	when  (format = 103 and rotate = 6) else
( "000000000000000000","000000011010010011","000000010001001010","000000010100001010","000000011010010011","000000000000000000")	when  (format = 103 and rotate = 7) else
( "000000000000000000","000000000000000000","011010010011000000","010001100010011000","011010001001010000","000011010010011000")	when  (format = 104 and rotate = 0) else
( "000000000000000000","000000000000000000","000000011010010011","000011010100001010","000010001001010011","000011010010011000")	when  (format = 104 and rotate = 1) else
( "000011010010011000","011010001001010000","010001100010011000","011010010011000000","000000000000000000","000000000000000000")	when  (format = 104 and rotate = 2) else
( "000011010010011000","000010001001010011","000011010100001010","000000011010010011","000000000000000000","000000000000000000")	when  (format = 104 and rotate = 3) else
( "000011010011000000","011010001010000000","010001100010000000","010001010011000000","011010011000000000","000000000000000000")	when  (format = 104 and rotate = 4) else
( "000000011010011000","000000010001010011","000000010100001010","000000011010001010","000000000011010011","000000000000000000")	when  (format = 104 and rotate = 5) else
( "000000000000000000","011010011000000000","010001010011000000","010001100010000000","011010001010000000","000011010011000000")	when  (format = 104 and rotate = 6) else
( "000000000000000000","000000000011010011","000000011010001010","000000010100001010","000000010001010011","000000011010011000")	when  (format = 104 and rotate = 7) else
( "000011010011000000","000010001010000000","011010001010000000","010001100010000000","010001010011000000","011010011000000000")	when  (format = 105 and rotate = 0) else
( "000000011010011000","000000010001010000","000000010001010011","000000010100001010","000000011010001010","000000000011010011")	when  (format = 105 and rotate = 1) else
( "011010011000000000","010001010011000000","010001100010000000","011010001010000000","000010001010000000","000011010011000000")	when  (format = 105 and rotate = 2) else
( "000000000011010011","000000011010001010","000000010100001010","000000010001010011","000000010001010000","000000011010011000")	when  (format = 105 and rotate = 3) else
( "011010010011000000","010001001010010011","011010100001001010","000011010010010011","000000000000000000","000000000000000000")	when  (format = 105 and rotate = 4) else
( "000000011010010011","011010010001001010","010001001100010011","011010010010011000","000000000000000000","000000000000000000")	when  (format = 105 and rotate = 5) else
( "000000000000000000","000000000000000000","000011010010010011","011010100001001010","010001001010010011","011010010011000000")	when  (format = 105 and rotate = 6) else
( "000000000000000000","000000000000000000","011010010010011000","010001001100010011","011010010001001010","000000011010010011")	when  (format = 105 and rotate = 7) else
( "000000000000000000","000011010011000000","011010001010000000","010001100010000000","010001001010000000","011010010011000000")	when  (format = 106 and rotate = 0) else
( "000000000000000000","000000011010011000","000000010001010011","000000010100001010","000000010001001010","000000011010010011")	when  (format = 106 and rotate = 1) else
( "011010010011000000","010001001010000000","010001100010000000","011010001010000000","000011010011000000","000000000000000000")	when  (format = 106 and rotate = 2) else
( "000000011010010011","000000010001001010","000000010100001010","000000010001010011","000000011010011000","000000000000000000")	when  (format = 106 and rotate = 3) else
( "011010010011000000","010001001010011000","010001100001010000","011010010010011000","000000000000000000","000000000000000000")	when  (format = 106 and rotate = 4) else
( "000000011010010011","000011010001001010","000010001100001010","000011010010010011","000000000000000000","000000000000000000")	when  (format = 106 and rotate = 5) else
( "000000000000000000","000000000000000000","011010010010011000","010001100001010000","010001001010011000","011010010011000000")	when  (format = 106 and rotate = 6) else
( "000000000000000000","000000000000000000","000011010010010011","000010001100001010","000011010001001010","000000011010010011")	when  (format = 106 and rotate = 7) else
( "000000000000000000","011010010011000000","010001001010000000","011010100010000000","010001001010000000","011010010011000000")	when  (format = 107 and rotate = 0) else
( "000000000000000000","000000011010010011","000000010001001010","000000010100010011","000000010001001010","000000011010010011")	when  (format = 107 and rotate = 1) else
( "011010010011000000","010001001010000000","011010100010000000","010001001010000000","011010010011000000","000000000000000000")	when  (format = 107 and rotate = 2) else
( "000000011010010011","000000010001001010","000000010100010011","000000010001001010","000000011010010011","000000000000000000")	when  (format = 107 and rotate = 3) else
( "011010011010011000","010001010001010000","010001100001010000","011010010010011000","000000000000000000","000000000000000000")	when  (format = 107 and rotate = 4) else
( "000011010011010011","000010001010001010","000010001100001010","000011010010010011","000000000000000000","000000000000000000")	when  (format = 107 and rotate = 5) else
( "000000000000000000","000000000000000000","011010010010011000","010001100001010000","010001010001010000","011010011010011000")	when  (format = 107 and rotate = 6) else
( "000000000000000000","000000000000000000","000011010010010011","000010001100001010","000010001010001010","000011010011010011")	when  (format = 107 and rotate = 7) else
( "000000000000000000","000011010011000000","000010001010000000","011010100010011000","010001001001010000","011010010010011000")	when  (format = 108 and rotate = 0) else
( "000000000000000000","000000011010011000","000000010001010000","000011010100010011","000010001001001010","000011010010010011")	when  (format = 108 and rotate = 1) else
( "011010010010011000","010001001001010000","011010100010011000","000010001010000000","000011010011000000","000000000000000000")	when  (format = 108 and rotate = 2) else
( "000011010010010011","000010001001001010","000011010100010011","000000010001010000","000000011010011000","000000000000000000")	when  (format = 108 and rotate = 3) else
( "011010011000000000","010001010010011000","010001100001010000","010001010010011000","011010011000000000","000000000000000000")	when  (format = 108 and rotate = 4) else
( "000000000011010011","000011010010001010","000010001100001010","000011010010001010","000000000011010011","000000000000000000")	when  (format = 108 and rotate = 5) else
( "000000000000000000","011010011000000000","010001010010011000","010001100001010000","010001010010011000","011010011000000000")	when  (format = 108 and rotate = 6) else
( "000000000000000000","000000000011010011","000011010010001010","000010001100001010","000011010010001010","000000000011010011")	when  (format = 108 and rotate = 7) else
( "000011010011000000","000010001010000000","000010001010010011","000010100001001010","000011010010010011","000000000000000000")	when  (format = 109 and rotate = 0) else
( "000000011010011000","000000010001010000","011010010001010000","010001001100010000","011010010010011000","000000000000000000")	when  (format = 109 and rotate = 1) else
( "000000000000000000","000011010010010011","000010100001001010","000010001010010011","000010001010000000","000011010011000000")	when  (format = 109 and rotate = 2) else
( "000000000000000000","011010010010011000","010001001100010000","011010010001010000","000000010001010000","000000011010011000")	when  (format = 109 and rotate = 3) else
( "000000000000000000","000011010010010011","000010100001001010","000010001010010011","000010001010000000","000011010011000000")	when  (format = 109 and rotate = 4) else
( "000000000000000000","011010010010011000","010001001100010000","011010010001010000","000000010001010000","000000011010011000")	when  (format = 109 and rotate = 5) else
( "000011010011000000","000010001010000000","000010001010010011","000010100001001010","000011010010010011","000000000000000000")	when  (format = 109 and rotate = 6) else
( "000000011010011000","000000010001010000","011010010001010000","010001001100010000","011010010010011000","000000000000000000")	when  (format = 109 and rotate = 7) else
( "000000000000000000","011010010011000000","010001001010011000","011010100001010000","000011010001010000","000000011010011000")	when  (format = 110 and rotate = 0) else
( "000000000000000000","000000011010010011","000011010001001010","000010001100010011","000010001010011000","000011010011000000")	when  (format = 110 and rotate = 1) else
( "000000011010011000","000011010001010000","011010100001010000","010001001010011000","011010010011000000","000000000000000000")	when  (format = 110 and rotate = 2) else
( "000011010011000000","000010001010011000","000010001100010011","000011010001001010","000000011010010011","000000000000000000")	when  (format = 110 and rotate = 3) else
( "000000011010011000","000011010001010000","011010100001010000","010001001010011000","011010010011000000","000000000000000000")	when  (format = 110 and rotate = 4) else
( "000011010011000000","000010001010011000","000010001100010011","000011010001001010","000000011010010011","000000000000000000")	when  (format = 110 and rotate = 5) else
( "000000000000000000","011010010011000000","010001001010011000","011010100001010000","000011010001010000","000000011010011000")	when  (format = 110 and rotate = 6) else
( "000000000000000000","000000011010010011","000011010001001010","000010001100010011","000010001010011000","000011010011000000")	when  (format = 110 and rotate = 7) else
( "000000000000000000","011010011000000000","010001010010011000","010001100001010000","011010010001010000","000000011010011000")	when  (format = 111 and rotate = 0) else
( "000000000000000000","000000000011010011","000011010010001010","000010001100001010","000010001010010011","000011010011000000")	when  (format = 111 and rotate = 1) else
( "000000011010011000","011010010001010000","010001100001010000","010001010010011000","011010011000000000","000000000000000000")	when  (format = 111 and rotate = 2) else
( "000011010011000000","000010001010010011","000010001100001010","000011010010001010","000000000011010011","000000000000000000")	when  (format = 111 and rotate = 3) else
( "000011010010011000","000010001001010000","011010100010011000","010001001010000000","011010010011000000","000000000000000000")	when  (format = 111 and rotate = 4) else
( "000011010010011000","000010001001010000","000011010100010011","000000010001001010","000000011010010011","000000000000000000")	when  (format = 111 and rotate = 5) else
( "000000000000000000","011010010011000000","010001001010000000","011010100010011000","000010001001010000","000011010010011000")	when  (format = 111 and rotate = 6) else
( "000000000000000000","000000011010010011","000000010001001010","000011010100010011","000010001001010000","000011010010011000")	when  (format = 111 and rotate = 7) else
( "000000000000000000","011010011000000000","010001010010011000","010001100001010000","011010001010011000","000011010011000000")	when  (format = 112 and rotate = 0) else
( "000000000000000000","000000000011010011","000011010010001010","000010001100001010","000011010001010011","000000011010011000")	when  (format = 112 and rotate = 1) else
( "000011010011000000","011010001010011000","010001100001010000","010001010010011000","011010011000000000","000000000000000000")	when  (format = 112 and rotate = 2) else
( "000000011010011000","000011010001010011","000010001100001010","000011010010001010","000000000011010011","000000000000000000")	when  (format = 112 and rotate = 3) else
( "000011010010011000","011010001001010000","010001100010011000","011010001010000000","000011010011000000","000000000000000000")	when  (format = 112 and rotate = 4) else
( "000011010010011000","000010001001010011","000011010100001010","000000010001010011","000000011010011000","000000000000000000")	when  (format = 112 and rotate = 5) else
( "000000000000000000","000011010011000000","011010001010000000","010001100010011000","011010001001010000","000011010010011000")	when  (format = 112 and rotate = 6) else
( "000000000000000000","000000011010011000","000000010001010011","000011010100001010","000010001001010011","000011010010011000")	when  (format = 112 and rotate = 7) else
( "000000000000000000","000011010011000000","011010001010011000","010001100001010000","011010001010011000","000011010011000000")	when  (format = 113 and rotate = 0) else
( "000000000000000000","000000011010011000","000011010001010011","000010001100001010","000011010001010011","000000011010011000")	when  (format = 113 and rotate = 1) else
( "000011010011000000","011010001010011000","010001100001010000","011010001010011000","000011010011000000","000000000000000000")	when  (format = 113 and rotate = 2) else
( "000000011010011000","000011010001010011","000010001100001010","000011010001010011","000000011010011000","000000000000000000")	when  (format = 113 and rotate = 3) else
( "000011010011000000","011010001010011000","010001100001010000","011010001010011000","000011010011000000","000000000000000000")	when  (format = 113 and rotate = 4) else
( "000000011010011000","000011010001010011","000010001100001010","000011010001010011","000000011010011000","000000000000000000")	when  (format = 113 and rotate = 5) else
( "000000000000000000","000011010011000000","011010001010011000","010001100001010000","011010001010011000","000011010011000000")	when  (format = 113 and rotate = 6) else
( "000000000000000000","000000011010011000","000011010001010011","000010001100001010","000011010001010011","000000011010011000") ;--	when  (format = 17 and rotate = 7) ;




data_decoded <= std_logic_vector(X_ini(4 downto 0)) & std_logic_vector(Y_ini(4 downto 0)) & sampler(5) & sampler(4) & sampler(3) & sampler(2) & sampler(1) & sampler(0);



	min_max_out <= mix_array(16) when (format = 97) else
						mix_array(15) when (format = 98) else
						mix_array(14) when (format = 99) else
						mix_array(13) when (format = 100) else
						mix_array(12) when (format = 101) else
						mix_array(11) when (format = 102) else
						mix_array(10) when (format = 103) else
						mix_array(9) when (format = 104) else
						mix_array(8) when (format = 105) else
						mix_array(7) when (format = 106) else
						mix_array(6) when (format = 107) else
						mix_array(5) when (format = 108) else
						mix_array(4) when (format = 109) else	
						mix_array(3) when (format = 110) else
						mix_array(2) when (format = 111) else
						mix_array(1) when (format = 112) else
						mix_array(0);

		alaki <= 

end Gate_level;


---------------------------------------------------------------------------------------------------------------------------------
architecture test_bench of program is

  -- Component Declaration
Component x Port ( datain : in std_logic_vector(31 downto 0);
				  data_decoded : out std_logic_vector (117 downto 0)
				  );
end component;
for g:x use Entity work.program(Gate_level);

signal datain1 : std_logic_vector(31 downto 0);
signal data_decoded1 : std_logic_vector (117 downto 0);
begin

-- Component Instantiation
  g: x PORT MAP(datain1,data_decoded1);
		 
    datain1 <= "01100001001101010110001000110110"; --"1100000000000000" after 2 ns,"1010101010101010" after 4 ns,"1111111111111111" after 6 ns,"1111111100000000" after 8 ns,"1111110011001001" after 10 ns; '1','0' after 10 ns;

end test_bench;



